-- Projekt Logikanalysator an der FH-Augsburg
-- 5. Semester, Technische Informatik,  WS2013/2014
-- A. Gareis, S. Vockinger
-- CPLD Komponente: eval_top_level für Einsatz auf dem TPLE-Board
-- Datum: 19.12.2013
-- Vers.: 1.0
-- ===========================================================================

library ieee;
use ieee.std_logic_1164.all;

entity top_level_tple is
	port (
		clk : in std_ulogic;
		ext_reset : in std_ulogic;
		
		-- mega Interface
		M_clk	: in std_ulogic;
		M_rw : in std_ulogic;
		M_nib_sel : in std_ulogic;
		M_reg_sel : in std_ulogic_vector(1 downto 0);
		M_data : inout std_logic_vector(3 downto 0);
		M_int : out std_ulogic;
		
		-- RAM Interface
		ram_data : inout std_logic_vector(15 downto 0);
		ram_adr : out std_ulogic_vector(17 downto 0);
		lb : out std_ulogic;
		ub : out std_ulogic;
		we : out std_ulogic;
		ce1 : out std_ulogic;
		ce2 : out std_ulogic;
		oe : out std_ulogic;
		
		-- Measure Interface
		io_dir : out std_ulogic;
		io_data : in std_ulogic_vector(23 downto 0)	--TODO: Change to : inout std_logic_vector(23 downto 0) when signals should be generated by tple
	);
end entity;

architecture structure of top_level_tple is

	component top_level
		port (
			clk : in std_ulogic;
			ext_reset : in std_ulogic;
			
			-- mega Interface
			M_clk	: in std_ulogic;
			M_rw : in std_ulogic;
			M_nib_sel : in std_ulogic;
			M_reg_sel : in std_ulogic_vector(1 downto 0);
			M_data : inout std_logic_vector(3 downto 0);
			M_int : out std_ulogic;
			
			--RAM Interface
			ram_data : inout std_logic_vector(15 downto 0);
			ram_adr : out std_ulogic_vector(17 downto 0);
			lb : out std_ulogic;
			ub : out std_ulogic;
			we : out std_ulogic;
			ce1 : out std_ulogic;
			ce2 : out std_ulogic;
			oe : out std_ulogic;
			
			-- Measure Interface
			io_dir : out std_ulogic;
			io_data : in std_ulogic_vector(7 downto 0)	--TODO: Change to : inout std_logic_vector(7 downto 0) when signals should be generated by tple
		);
	end component;

	signal used_io_pins : std_ulogic_vector(7 downto 0);
	
begin

	used_io_pins <=  io_data(23 downto 20) & io_data(3 downto 0);
	
	topLevel : top_level
		port map (
			clk => clk,
			ext_reset => ext_reset,
			-- mega Interface
			M_clk	=> M_clk,
			M_rw => M_rw,
			M_nib_sel => M_nib_sel,
			M_reg_sel => M_reg_sel,
			M_data => M_data,
			M_int => M_int,
			--RAM Interface
			ram_data => ram_data,
			ram_adr => ram_adr,
			lb => lb,
			ub => ub,
			we => we,
			ce1 => ce1,
			ce2 => ce2,
			oe => oe,
			io_dir => io_dir,
			io_data => used_io_pins 
		);

end architecture;