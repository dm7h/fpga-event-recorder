-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2015.04.27409

-- Build Date:         May 27 2015 16:13:32

-- File Generated:     Feb 6 2017 16:52:13

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "gpio_pwm" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of gpio_pwm
entity gpio_pwm is
port (
    pwm_prescale : in std_logic_vector(2 downto 0);
    pwm_ctrl : in std_logic_vector(1 downto 0);
    pwm_hout : in std_logic_vector(11 downto 0);
    pwm_lout : in std_logic_vector(11 downto 0);
    clk : in std_logic;
    pwm_pin : out std_logic;
    reset : in std_logic);
end gpio_pwm;

-- Architecture of gpio_pwm
-- View name is \INTERFACE\
architecture \INTERFACE\ of gpio_pwm is

signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4599\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4596\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4593\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3936\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3775\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3729\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3654\ : std_logic;
signal \N__3651\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3576\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3564\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3549\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3519\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3513\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3477\ : std_logic;
signal \N__3474\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3468\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3441\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3381\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3321\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3228\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3192\ : std_logic;
signal \N__3189\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3021\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2990\ : std_logic;
signal \N__2987\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2947\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2922\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2884\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2704\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2533\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2494\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2392\ : std_logic;
signal \N__2389\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2374\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2359\ : std_logic;
signal \N__2356\ : std_logic;
signal \N__2353\ : std_logic;
signal \N__2350\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2332\ : std_logic;
signal \N__2329\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \N__2317\ : std_logic;
signal \N__2314\ : std_logic;
signal \N__2311\ : std_logic;
signal \N__2308\ : std_logic;
signal \N__2305\ : std_logic;
signal \N__2302\ : std_logic;
signal \N__2299\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2287\ : std_logic;
signal \N__2284\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2275\ : std_logic;
signal \N__2272\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal pwm_pin_c : std_logic;
signal pwm_lout_c_9 : std_logic;
signal pwm_lout_c_6 : std_logic;
signal pwm_hout_c_9 : std_logic;
signal pwm_hout_c_8 : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal proc_pwm_fsm_pwm_loc8_0_data_tmp_0 : std_logic;
signal proc_pwm_fsm_pwm_loc8_0_data_tmp_1 : std_logic;
signal proc_pwm_fsm_pwm_loc8_0_data_tmp_2 : std_logic;
signal proc_pwm_fsm_pwm_loc8_0_data_tmp_3 : std_logic;
signal proc_pwm_fsm_pwm_loc8_0_data_tmp_4 : std_logic;
signal proc_pwm_fsm_pwm_loc8 : std_logic;
signal \pwm_lout_p1Z0Z_6\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_26\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_6\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_16\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_21\ : std_logic;
signal \pwm_hout_p1Z0Z_8\ : std_logic;
signal \pwm_hout_p1Z0Z_9\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_11\ : std_logic;
signal pwm_hout_c_5 : std_logic;
signal \pwm_hout_p1Z0Z_5\ : std_logic;
signal pwm_hout_c_4 : std_logic;
signal \pwm_hout_p1Z0Z_4\ : std_logic;
signal pwm_hout_c_0 : std_logic;
signal \pwm_hout_p1Z0Z_0\ : std_logic;
signal pwm_hout_c_3 : std_logic;
signal \pwm_hout_p1Z0Z_3\ : std_logic;
signal pwm_lout_c_2 : std_logic;
signal \pwm_lout_p1Z0Z_2\ : std_logic;
signal pwm_hout_c_1 : std_logic;
signal \pwm_hout_p1Z0Z_1\ : std_logic;
signal pwm_hout_c_2 : std_logic;
signal \pwm_hout_p1Z0Z_2\ : std_logic;
signal pwm_lout_c_3 : std_logic;
signal \pwm_lout_p1Z0Z_3\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_0_N_1\ : std_logic;
signal pwm_hout_c_6 : std_logic;
signal \pwm_hout_p1Z0Z_6\ : std_logic;
signal pwm_hout_c_10 : std_logic;
signal \pwm_hout_p1Z0Z_10\ : std_logic;
signal pwm_hout_c_7 : std_logic;
signal \pwm_hout_p1Z0Z_7\ : std_logic;
signal pwm_hout_c_11 : std_logic;
signal \pwm_hout_p1Z0Z_11\ : std_logic;
signal pwm_prescale_c_0 : std_logic;
signal pwm_lout_c_7 : std_logic;
signal \pwm_lout_p1Z0Z_7\ : std_logic;
signal pwm_prescale_c_2 : std_logic;
signal pwm_lout_c_8 : std_logic;
signal pwm_ctrl_c_0 : std_logic;
signal \pwm_lout_p1Z0Z_8\ : std_logic;
signal \pwm_lout_p1Z0Z_9\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_21\ : std_logic;
signal proc_pwm_fsm_pwm_loc20_0_data_tmp_0 : std_logic;
signal proc_pwm_fsm_pwm_loc20_0_data_tmp_1 : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_6\ : std_logic;
signal proc_pwm_fsm_pwm_loc20_0_data_tmp_2 : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_11\ : std_logic;
signal proc_pwm_fsm_pwm_loc20_0_data_tmp_3 : std_logic;
signal proc_pwm_fsm_pwm_loc20_0_data_tmp_4 : std_logic;
signal proc_pwm_fsm_pwm_loc20 : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal pwm_cnt_cry_0 : std_logic;
signal \pwm_cntZ0Z_2\ : std_logic;
signal pwm_cnt_cry_1 : std_logic;
signal \pwm_cntZ0Z_3\ : std_logic;
signal pwm_cnt_cry_2 : std_logic;
signal pwm_cnt_cry_3 : std_logic;
signal pwm_cnt_cry_4 : std_logic;
signal \pwm_cntZ0Z_6\ : std_logic;
signal pwm_cnt_cry_5 : std_logic;
signal \pwm_cntZ0Z_7\ : std_logic;
signal pwm_cnt_cry_6 : std_logic;
signal pwm_cnt_cry_7 : std_logic;
signal \pwm_cntZ0Z_8\ : std_logic;
signal \bfn_2_12_0_\ : std_logic;
signal \pwm_cntZ0Z_9\ : std_logic;
signal pwm_cnt_cry_8 : std_logic;
signal pwm_cnt_cry_9 : std_logic;
signal pwm_cnt_cry_10 : std_logic;
signal \N_8_cascade_\ : std_logic;
signal \prescale_cnt_p1Z0Z_0\ : std_logic;
signal \prescale_cnt_p1Z0Z_1\ : std_logic;
signal \N_38\ : std_logic;
signal \pwm_cntZ0Z_11\ : std_logic;
signal \pwm_cntZ0Z_10\ : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_1\ : std_logic;
signal pwm_lout_c_11 : std_logic;
signal \pwm_lout_p1Z0Z_11\ : std_logic;
signal pwm_lout_c_10 : std_logic;
signal \pwm_lout_p1Z0Z_10\ : std_logic;
signal pwm_lout_c_1 : std_logic;
signal pwm_ctrl_c_1 : std_logic;
signal pwm_lout_c_0 : std_logic;
signal \prescale_stop_p1Z0Z_6\ : std_logic;
signal \prescale_cnt_p1Z0Z_7\ : std_logic;
signal \prescale_stop_p1Z0Z_7\ : std_logic;
signal \prescale_cnt_p1Z0Z_6\ : std_logic;
signal \prescale_stop_p1Z0Z_10\ : std_logic;
signal \prescale_cnt_p1Z0Z_11\ : std_logic;
signal \prescale_cnt_p1Z0Z_10\ : std_logic;
signal \pwm_cntZ0Z_1\ : std_logic;
signal \pwm_lout_p1Z0Z_1\ : std_logic;
signal \pwm_cntZ0Z_0\ : std_logic;
signal \pwm_lout_p1Z0Z_0\ : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_26\ : std_logic;
signal \pwm_cntZ0Z_5\ : std_logic;
signal \pwm_cntZ0Z_4\ : std_logic;
signal \proc_pwm_fsm_pwm_loc20_0_N_16\ : std_logic;
signal \pwm_ctrl_p1Z0Z_0\ : std_logic;
signal \pwm_ctrl_p1Z0Z_1\ : std_logic;
signal \pwm_loc_1_sqmuxa_cascade_\ : std_logic;
signal \un1_pwm_loc8_1_0_cascade_\ : std_logic;
signal pwm_cnte_0_i : std_logic;
signal un1_pwm_loc8_1_0 : std_logic;
signal \prescale_tickZ0\ : std_logic;
signal pwm_loc_1_sqmuxa : std_logic;
signal pwm_loc_0_sqmuxa_1 : std_logic;
signal \pwm_loc_1_sqmuxa_1_cascade_\ : std_logic;
signal \pwm_locZ0\ : std_logic;
signal \proc_pwm_fsm_pwm_loc20_THRU_CO\ : std_logic;
signal \N_87\ : std_logic;
signal \pwm_toglZ0\ : std_logic;
signal \N_86\ : std_logic;
signal \N_87_cascade_\ : std_logic;
signal \proc_pwm_fsm_pwm_loc8_THRU_CO\ : std_logic;
signal \N_78_0_i\ : std_logic;
signal \prescale_cntZ0Z_0\ : std_logic;
signal prescale_cnt_s_0 : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \prescale_cntZ0Z_1\ : std_logic;
signal prescale_cnt_cry_0 : std_logic;
signal prescale_cnt_cry_1 : std_logic;
signal prescale_cnt_cry_2 : std_logic;
signal prescale_cnt_cry_3 : std_logic;
signal prescale_cnt_cry_4 : std_logic;
signal \prescale_cntZ0Z_6\ : std_logic;
signal prescale_cnt_cry_5 : std_logic;
signal \prescale_cntZ0Z_7\ : std_logic;
signal prescale_cnt_cry_6 : std_logic;
signal prescale_cnt_cry_7 : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal prescale_cnt_cry_8 : std_logic;
signal \prescale_cntZ0Z_10\ : std_logic;
signal prescale_cnt_cry_9 : std_logic;
signal \prescale_cntZ0Z_11\ : std_logic;
signal prescale_cnt_cry_10 : std_logic;
signal prescale_cnt_cry_11 : std_logic;
signal prescale_cnt_cry_12 : std_logic;
signal prescale_cnt_cry_13 : std_logic;
signal prescale_cnt_cry_14 : std_logic;
signal prescale_cnt_cry_15 : std_logic;
signal \N_8\ : std_logic;
signal \bfn_3_14_0_\ : std_logic;
signal \prescale_stop_p1Z0Z_0\ : std_logic;
signal \prescale_stop_p1Z0Z_1\ : std_logic;
signal pwm_lout_c_4 : std_logic;
signal \pwm_lout_p1Z0Z_4\ : std_logic;
signal \prescale_cntZ0Z_5\ : std_logic;
signal \prescale_stop_p1Z0Z_15\ : std_logic;
signal \prescale_cntZ0Z_14\ : std_logic;
signal \prescale_cnt_p1Z0Z_14\ : std_logic;
signal \prescale_cntZ0Z_15\ : std_logic;
signal \prescale_cnt_p1Z0Z_15\ : std_logic;
signal pwm_prescale_c_1 : std_logic;
signal pwm_lout_c_5 : std_logic;
signal \pwm_lout_p1Z0Z_5\ : std_logic;
signal \prescale_stop_p1Z0Z_8\ : std_logic;
signal \prescale_cntZ0Z_8\ : std_logic;
signal \prescale_cnt_p1Z0Z_8\ : std_logic;
signal \prescale_cntZ0Z_9\ : std_logic;
signal \prescale_cnt_p1Z0Z_9\ : std_logic;
signal \prescale_stop_p1Z0Z_2\ : std_logic;
signal \prescale_stop_p1Z0Z_3\ : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_41\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_1\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_0 : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_1 : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_11\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_2 : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_16\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_3 : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_21\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_4 : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_5 : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_31\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_6 : std_logic;
signal proc_pwm_cnt_prescale_cnt10_0_data_tmp_7 : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal proc_pwm_cnt_prescale_cnt10 : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_THRU_CO\ : std_logic;
signal \prescale_cnt_p1Z0Z_5\ : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_6\ : std_logic;
signal \prescale_stop_p1Z0Z_14\ : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_36\ : std_logic;
signal \prescale_cntZ0Z_12\ : std_logic;
signal \prescale_cntZ0Z_16\ : std_logic;
signal \prescale_cnt_p1Z0Z_16\ : std_logic;
signal \prescale_stop_p1Z0Z_5\ : std_logic;
signal prescale_stop_1_7 : std_logic;
signal \prescale_cntZ0Z_3\ : std_logic;
signal \prescale_cnt_p1Z0Z_3\ : std_logic;
signal \prescale_cntZ0Z_2\ : std_logic;
signal \prescale_cnt_p1Z0Z_2\ : std_logic;
signal \prescale_cntZ0Z_13\ : std_logic;
signal \prescale_stop_p1Z0Z_4\ : std_logic;
signal \prescale_cntZ0Z_4\ : std_logic;
signal \prescale_cnt_p1Z0Z_4\ : std_logic;
signal \pwm_prescale_p1Z0Z_2\ : std_logic;
signal \pwm_prescale_p1Z0Z_1\ : std_logic;
signal \prescale_cnt_p1Z0Z_13\ : std_logic;
signal \prescale_cnt_p1Z0Z_12\ : std_logic;
signal \proc_pwm_cnt_prescale_cnt10_0_N_26\ : std_logic;
signal prescale_stop_1_8 : std_logic;
signal \pwm_prescale_p1Z0Z_0\ : std_logic;
signal \prescale_stop_p1Z0Z_13\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_c_g : std_logic;
signal reset_c_g : std_logic;

signal reset_wire : std_logic;
signal clk_wire : std_logic;
signal pwm_hout_wire : std_logic_vector(11 downto 0);
signal pwm_lout_wire : std_logic_vector(11 downto 0);
signal pwm_ctrl_wire : std_logic_vector(1 downto 0);
signal pwm_prescale_wire : std_logic_vector(2 downto 0);
signal pwm_pin_wire : std_logic;

begin
    reset_wire <= reset;
    clk_wire <= clk;
    pwm_hout_wire <= pwm_hout;
    pwm_lout_wire <= pwm_lout;
    pwm_ctrl_wire <= pwm_ctrl;
    pwm_prescale_wire <= pwm_prescale;
    pwm_pin <= pwm_pin_wire;

    \reset_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5028\,
            GLOBALBUFFEROUTPUT => reset_c_g
        );

    \reset_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5030\,
            DIN => \N__5029\,
            DOUT => \N__5028\,
            PACKAGEPIN => reset_wire
        );

    \reset_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5030\,
            PADOUT => \N__5029\,
            PADIN => \N__5028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__5018\,
            GLOBALBUFFEROUTPUT => clk_c_g
        );

    \clk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5020\,
            DIN => \N__5019\,
            DOUT => \N__5018\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5020\,
            PADOUT => \N__5019\,
            PADIN => \N__5018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5009\,
            DIN => \N__5008\,
            DOUT => \N__5007\,
            PACKAGEPIN => pwm_hout_wire(11)
        );

    \pwm_hout_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5009\,
            PADOUT => \N__5008\,
            PADIN => \N__5007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_11,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__5000\,
            DIN => \N__4999\,
            DOUT => \N__4998\,
            PACKAGEPIN => pwm_hout_wire(5)
        );

    \pwm_hout_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__5000\,
            PADOUT => \N__4999\,
            PADIN => \N__4998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4991\,
            DIN => \N__4990\,
            DOUT => \N__4989\,
            PACKAGEPIN => pwm_hout_wire(2)
        );

    \pwm_hout_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4991\,
            PADOUT => \N__4990\,
            PADIN => \N__4989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4982\,
            DIN => \N__4981\,
            DOUT => \N__4980\,
            PACKAGEPIN => pwm_lout_wire(4)
        );

    \pwm_lout_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4982\,
            PADOUT => \N__4981\,
            PADIN => \N__4980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_ctrl_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4973\,
            DIN => \N__4972\,
            DOUT => \N__4971\,
            PACKAGEPIN => pwm_ctrl_wire(0)
        );

    \pwm_ctrl_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4973\,
            PADOUT => \N__4972\,
            PADIN => \N__4971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_ctrl_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4964\,
            DIN => \N__4963\,
            DOUT => \N__4962\,
            PACKAGEPIN => pwm_lout_wire(9)
        );

    \pwm_lout_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4964\,
            PADOUT => \N__4963\,
            PADIN => \N__4962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_9,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_prescale_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4955\,
            DIN => \N__4954\,
            DOUT => \N__4953\,
            PACKAGEPIN => pwm_prescale_wire(1)
        );

    \pwm_prescale_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4955\,
            PADOUT => \N__4954\,
            PADIN => \N__4953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_prescale_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4946\,
            DIN => \N__4945\,
            DOUT => \N__4944\,
            PACKAGEPIN => pwm_hout_wire(7)
        );

    \pwm_hout_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4946\,
            PADOUT => \N__4945\,
            PADIN => \N__4944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4937\,
            DIN => \N__4936\,
            DOUT => \N__4935\,
            PACKAGEPIN => pwm_lout_wire(1)
        );

    \pwm_lout_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4937\,
            PADOUT => \N__4936\,
            PADIN => \N__4935\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_pin_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4928\,
            DIN => \N__4927\,
            DOUT => \N__4926\,
            PACKAGEPIN => pwm_pin_wire
        );

    \pwm_pin_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__4928\,
            PADOUT => \N__4927\,
            PADIN => \N__4926\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4919\,
            DIN => \N__4918\,
            DOUT => \N__4917\,
            PACKAGEPIN => pwm_lout_wire(6)
        );

    \pwm_lout_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4919\,
            PADOUT => \N__4918\,
            PADIN => \N__4917\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4910\,
            DIN => \N__4909\,
            DOUT => \N__4908\,
            PACKAGEPIN => pwm_hout_wire(9)
        );

    \pwm_hout_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4910\,
            PADOUT => \N__4909\,
            PADIN => \N__4908\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_9,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4901\,
            DIN => \N__4900\,
            DOUT => \N__4899\,
            PACKAGEPIN => pwm_hout_wire(4)
        );

    \pwm_hout_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4901\,
            PADOUT => \N__4900\,
            PADIN => \N__4899\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4892\,
            DIN => \N__4891\,
            DOUT => \N__4890\,
            PACKAGEPIN => pwm_hout_wire(1)
        );

    \pwm_hout_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4892\,
            PADOUT => \N__4891\,
            PADIN => \N__4890\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4883\,
            DIN => \N__4882\,
            DOUT => \N__4881\,
            PACKAGEPIN => pwm_lout_wire(3)
        );

    \pwm_lout_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4883\,
            PADOUT => \N__4882\,
            PADIN => \N__4881\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_ctrl_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4874\,
            DIN => \N__4873\,
            DOUT => \N__4872\,
            PACKAGEPIN => pwm_ctrl_wire(1)
        );

    \pwm_ctrl_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4874\,
            PADOUT => \N__4873\,
            PADIN => \N__4872\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_ctrl_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_prescale_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4865\,
            DIN => \N__4864\,
            DOUT => \N__4863\,
            PACKAGEPIN => pwm_prescale_wire(2)
        );

    \pwm_prescale_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4865\,
            PADOUT => \N__4864\,
            PADIN => \N__4863\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_prescale_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4856\,
            DIN => \N__4855\,
            DOUT => \N__4854\,
            PACKAGEPIN => pwm_lout_wire(10)
        );

    \pwm_lout_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4856\,
            PADOUT => \N__4855\,
            PADIN => \N__4854\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_10,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4847\,
            DIN => \N__4846\,
            DOUT => \N__4845\,
            PACKAGEPIN => pwm_lout_wire(8)
        );

    \pwm_lout_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4847\,
            PADOUT => \N__4846\,
            PADIN => \N__4845\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_8,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4838\,
            DIN => \N__4837\,
            DOUT => \N__4836\,
            PACKAGEPIN => pwm_hout_wire(10)
        );

    \pwm_hout_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4838\,
            PADOUT => \N__4837\,
            PADIN => \N__4836\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_10,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4829\,
            DIN => \N__4828\,
            DOUT => \N__4827\,
            PACKAGEPIN => pwm_hout_wire(6)
        );

    \pwm_hout_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4829\,
            PADOUT => \N__4828\,
            PADIN => \N__4827\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4820\,
            DIN => \N__4819\,
            DOUT => \N__4818\,
            PACKAGEPIN => pwm_lout_wire(0)
        );

    \pwm_lout_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4820\,
            PADOUT => \N__4819\,
            PADIN => \N__4818\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4811\,
            DIN => \N__4810\,
            DOUT => \N__4809\,
            PACKAGEPIN => pwm_hout_wire(3)
        );

    \pwm_hout_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4811\,
            PADOUT => \N__4810\,
            PADIN => \N__4809\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4802\,
            DIN => \N__4801\,
            DOUT => \N__4800\,
            PACKAGEPIN => pwm_lout_wire(5)
        );

    \pwm_lout_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4802\,
            PADOUT => \N__4801\,
            PADIN => \N__4800\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4793\,
            DIN => \N__4792\,
            DOUT => \N__4791\,
            PACKAGEPIN => pwm_hout_wire(8)
        );

    \pwm_hout_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4793\,
            PADOUT => \N__4792\,
            PADIN => \N__4791\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_8,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_prescale_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4784\,
            DIN => \N__4783\,
            DOUT => \N__4782\,
            PACKAGEPIN => pwm_prescale_wire(0)
        );

    \pwm_prescale_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4784\,
            PADOUT => \N__4783\,
            PADIN => \N__4782\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_prescale_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_hout_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4775\,
            DIN => \N__4774\,
            DOUT => \N__4773\,
            PACKAGEPIN => pwm_hout_wire(0)
        );

    \pwm_hout_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4775\,
            PADOUT => \N__4774\,
            PADIN => \N__4773\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_hout_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4766\,
            DIN => \N__4765\,
            DOUT => \N__4764\,
            PACKAGEPIN => pwm_lout_wire(2)
        );

    \pwm_lout_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4766\,
            PADOUT => \N__4765\,
            PADIN => \N__4764\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4757\,
            DIN => \N__4756\,
            DOUT => \N__4755\,
            PACKAGEPIN => pwm_lout_wire(11)
        );

    \pwm_lout_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4757\,
            PADOUT => \N__4756\,
            PADIN => \N__4755\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_11,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pwm_lout_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4748\,
            DIN => \N__4747\,
            DOUT => \N__4746\,
            PACKAGEPIN => pwm_lout_wire(7)
        );

    \pwm_lout_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__4748\,
            PADOUT => \N__4747\,
            PADIN => \N__4746\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => pwm_lout_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1020\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4723\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4723\,
            I => \prescale_stop_p1Z0Z_4\
        );

    \I__1017\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4717\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__4717\,
            I => \N__4713\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4710\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__4713\,
            I => \prescale_cntZ0Z_4\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__4710\,
            I => \prescale_cntZ0Z_4\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4702\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4702\,
            I => \prescale_cnt_p1Z0Z_4\
        );

    \I__1010\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__1009\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4690\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4684\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4681\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4693\,
            I => \N__4673\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4690\,
            I => \N__4673\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4668\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4668\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4662\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4657\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4657\
        );

    \I__999\ : InMux
    port map (
            O => \N__4680\,
            I => \N__4654\
        );

    \I__998\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4649\
        );

    \I__997\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4649\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__4673\,
            I => \N__4643\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4643\
        );

    \I__994\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4636\
        );

    \I__993\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4636\
        );

    \I__992\ : InMux
    port map (
            O => \N__4665\,
            I => \N__4636\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4629\
        );

    \I__990\ : Span4Mux_v
    port map (
            O => \N__4657\,
            I => \N__4629\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__4654\,
            I => \N__4629\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__4649\,
            I => \N__4626\
        );

    \I__987\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4623\
        );

    \I__986\ : Span4Mux_h
    port map (
            O => \N__4643\,
            I => \N__4620\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4636\,
            I => \N__4615\
        );

    \I__984\ : Span4Mux_h
    port map (
            O => \N__4629\,
            I => \N__4615\
        );

    \I__983\ : Span12Mux_h
    port map (
            O => \N__4626\,
            I => \N__4610\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4623\,
            I => \N__4610\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__4620\,
            I => \pwm_prescale_p1Z0Z_2\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__4615\,
            I => \pwm_prescale_p1Z0Z_2\
        );

    \I__979\ : Odrv12
    port map (
            O => \N__4610\,
            I => \pwm_prescale_p1Z0Z_2\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__977\ : InMux
    port map (
            O => \N__4600\,
            I => \N__4588\
        );

    \I__976\ : InMux
    port map (
            O => \N__4599\,
            I => \N__4588\
        );

    \I__975\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4585\
        );

    \I__974\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4582\
        );

    \I__973\ : InMux
    port map (
            O => \N__4596\,
            I => \N__4579\
        );

    \I__972\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4576\
        );

    \I__971\ : InMux
    port map (
            O => \N__4594\,
            I => \N__4569\
        );

    \I__970\ : InMux
    port map (
            O => \N__4593\,
            I => \N__4566\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__4588\,
            I => \N__4563\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__4585\,
            I => \N__4556\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4582\,
            I => \N__4556\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4579\,
            I => \N__4556\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4576\,
            I => \N__4553\
        );

    \I__964\ : InMux
    port map (
            O => \N__4575\,
            I => \N__4550\
        );

    \I__963\ : InMux
    port map (
            O => \N__4574\,
            I => \N__4545\
        );

    \I__962\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4545\
        );

    \I__961\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4542\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4569\,
            I => \N__4537\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4566\,
            I => \N__4537\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__4563\,
            I => \N__4532\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__4556\,
            I => \N__4532\
        );

    \I__956\ : Odrv12
    port map (
            O => \N__4553\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4550\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__4545\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4542\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__4537\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__4532\,
            I => \pwm_prescale_p1Z0Z_1\
        );

    \I__950\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__4513\,
            I => \prescale_cnt_p1Z0Z_13\
        );

    \I__947\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4507\,
            I => \prescale_cnt_p1Z0Z_12\
        );

    \I__945\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4501\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_26\
        );

    \I__943\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4495\,
            I => prescale_stop_1_8
        );

    \I__941\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4481\
        );

    \I__940\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4481\
        );

    \I__939\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4481\
        );

    \I__938\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4475\
        );

    \I__937\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4472\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4481\,
            I => \N__4469\
        );

    \I__935\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4466\
        );

    \I__934\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4463\
        );

    \I__933\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4458\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4475\,
            I => \N__4453\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4472\,
            I => \N__4453\
        );

    \I__930\ : Span4Mux_v
    port map (
            O => \N__4469\,
            I => \N__4450\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4466\,
            I => \N__4445\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4463\,
            I => \N__4445\
        );

    \I__927\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4440\
        );

    \I__926\ : InMux
    port map (
            O => \N__4461\,
            I => \N__4440\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__4458\,
            I => \N__4435\
        );

    \I__924\ : Span4Mux_v
    port map (
            O => \N__4453\,
            I => \N__4435\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__4450\,
            I => \N__4427\
        );

    \I__922\ : Span4Mux_h
    port map (
            O => \N__4445\,
            I => \N__4427\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4440\,
            I => \N__4427\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__4435\,
            I => \N__4424\
        );

    \I__919\ : InMux
    port map (
            O => \N__4434\,
            I => \N__4421\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__4427\,
            I => \pwm_prescale_p1Z0Z_0\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__4424\,
            I => \pwm_prescale_p1Z0Z_0\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__4421\,
            I => \pwm_prescale_p1Z0Z_0\
        );

    \I__915\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__4411\,
            I => \prescale_stop_p1Z0Z_13\
        );

    \I__913\ : ClkMux
    port map (
            O => \N__4408\,
            I => \N__4333\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4407\,
            I => \N__4333\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4406\,
            I => \N__4333\
        );

    \I__910\ : ClkMux
    port map (
            O => \N__4405\,
            I => \N__4333\
        );

    \I__909\ : ClkMux
    port map (
            O => \N__4404\,
            I => \N__4333\
        );

    \I__908\ : ClkMux
    port map (
            O => \N__4403\,
            I => \N__4333\
        );

    \I__907\ : ClkMux
    port map (
            O => \N__4402\,
            I => \N__4333\
        );

    \I__906\ : ClkMux
    port map (
            O => \N__4401\,
            I => \N__4333\
        );

    \I__905\ : ClkMux
    port map (
            O => \N__4400\,
            I => \N__4333\
        );

    \I__904\ : ClkMux
    port map (
            O => \N__4399\,
            I => \N__4333\
        );

    \I__903\ : ClkMux
    port map (
            O => \N__4398\,
            I => \N__4333\
        );

    \I__902\ : ClkMux
    port map (
            O => \N__4397\,
            I => \N__4333\
        );

    \I__901\ : ClkMux
    port map (
            O => \N__4396\,
            I => \N__4333\
        );

    \I__900\ : ClkMux
    port map (
            O => \N__4395\,
            I => \N__4333\
        );

    \I__899\ : ClkMux
    port map (
            O => \N__4394\,
            I => \N__4333\
        );

    \I__898\ : ClkMux
    port map (
            O => \N__4393\,
            I => \N__4333\
        );

    \I__897\ : ClkMux
    port map (
            O => \N__4392\,
            I => \N__4333\
        );

    \I__896\ : ClkMux
    port map (
            O => \N__4391\,
            I => \N__4333\
        );

    \I__895\ : ClkMux
    port map (
            O => \N__4390\,
            I => \N__4333\
        );

    \I__894\ : ClkMux
    port map (
            O => \N__4389\,
            I => \N__4333\
        );

    \I__893\ : ClkMux
    port map (
            O => \N__4388\,
            I => \N__4333\
        );

    \I__892\ : ClkMux
    port map (
            O => \N__4387\,
            I => \N__4333\
        );

    \I__891\ : ClkMux
    port map (
            O => \N__4386\,
            I => \N__4333\
        );

    \I__890\ : ClkMux
    port map (
            O => \N__4385\,
            I => \N__4333\
        );

    \I__889\ : ClkMux
    port map (
            O => \N__4384\,
            I => \N__4333\
        );

    \I__888\ : GlobalMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__887\ : gio2CtrlBuf
    port map (
            O => \N__4330\,
            I => clk_c_g
        );

    \I__886\ : SRMux
    port map (
            O => \N__4327\,
            I => \N__4252\
        );

    \I__885\ : SRMux
    port map (
            O => \N__4326\,
            I => \N__4252\
        );

    \I__884\ : SRMux
    port map (
            O => \N__4325\,
            I => \N__4252\
        );

    \I__883\ : SRMux
    port map (
            O => \N__4324\,
            I => \N__4252\
        );

    \I__882\ : SRMux
    port map (
            O => \N__4323\,
            I => \N__4252\
        );

    \I__881\ : SRMux
    port map (
            O => \N__4322\,
            I => \N__4252\
        );

    \I__880\ : SRMux
    port map (
            O => \N__4321\,
            I => \N__4252\
        );

    \I__879\ : SRMux
    port map (
            O => \N__4320\,
            I => \N__4252\
        );

    \I__878\ : SRMux
    port map (
            O => \N__4319\,
            I => \N__4252\
        );

    \I__877\ : SRMux
    port map (
            O => \N__4318\,
            I => \N__4252\
        );

    \I__876\ : SRMux
    port map (
            O => \N__4317\,
            I => \N__4252\
        );

    \I__875\ : SRMux
    port map (
            O => \N__4316\,
            I => \N__4252\
        );

    \I__874\ : SRMux
    port map (
            O => \N__4315\,
            I => \N__4252\
        );

    \I__873\ : SRMux
    port map (
            O => \N__4314\,
            I => \N__4252\
        );

    \I__872\ : SRMux
    port map (
            O => \N__4313\,
            I => \N__4252\
        );

    \I__871\ : SRMux
    port map (
            O => \N__4312\,
            I => \N__4252\
        );

    \I__870\ : SRMux
    port map (
            O => \N__4311\,
            I => \N__4252\
        );

    \I__869\ : SRMux
    port map (
            O => \N__4310\,
            I => \N__4252\
        );

    \I__868\ : SRMux
    port map (
            O => \N__4309\,
            I => \N__4252\
        );

    \I__867\ : SRMux
    port map (
            O => \N__4308\,
            I => \N__4252\
        );

    \I__866\ : SRMux
    port map (
            O => \N__4307\,
            I => \N__4252\
        );

    \I__865\ : SRMux
    port map (
            O => \N__4306\,
            I => \N__4252\
        );

    \I__864\ : SRMux
    port map (
            O => \N__4305\,
            I => \N__4252\
        );

    \I__863\ : SRMux
    port map (
            O => \N__4304\,
            I => \N__4252\
        );

    \I__862\ : SRMux
    port map (
            O => \N__4303\,
            I => \N__4252\
        );

    \I__861\ : GlobalMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__860\ : gio2CtrlBuf
    port map (
            O => \N__4249\,
            I => reset_c_g
        );

    \I__859\ : InMux
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__4240\,
            I => \prescale_cnt_p1Z0Z_5\
        );

    \I__856\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4234\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_6\
        );

    \I__854\ : InMux
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4228\,
            I => \N__4224\
        );

    \I__852\ : InMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__851\ : Odrv12
    port map (
            O => \N__4224\,
            I => \prescale_stop_p1Z0Z_14\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4221\,
            I => \prescale_stop_p1Z0Z_14\
        );

    \I__849\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4213\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4213\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_36\
        );

    \I__847\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__4204\,
            I => \N__4200\
        );

    \I__844\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4197\
        );

    \I__843\ : Odrv4
    port map (
            O => \N__4200\,
            I => \prescale_cntZ0Z_12\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4197\,
            I => \prescale_cntZ0Z_12\
        );

    \I__841\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4189\,
            I => \N__4185\
        );

    \I__839\ : InMux
    port map (
            O => \N__4188\,
            I => \N__4182\
        );

    \I__838\ : Odrv4
    port map (
            O => \N__4185\,
            I => \prescale_cntZ0Z_16\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4182\,
            I => \prescale_cntZ0Z_16\
        );

    \I__836\ : InMux
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4174\,
            I => \prescale_cnt_p1Z0Z_16\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__833\ : InMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4165\,
            I => \prescale_stop_p1Z0Z_5\
        );

    \I__831\ : InMux
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4159\,
            I => prescale_stop_1_7
        );

    \I__829\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4150\,
            I => \N__4146\
        );

    \I__826\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4143\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__4146\,
            I => \prescale_cntZ0Z_3\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4143\,
            I => \prescale_cntZ0Z_3\
        );

    \I__823\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4135\,
            I => \prescale_cnt_p1Z0Z_3\
        );

    \I__821\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4129\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__819\ : Span4Mux_h
    port map (
            O => \N__4126\,
            I => \N__4122\
        );

    \I__818\ : InMux
    port map (
            O => \N__4125\,
            I => \N__4119\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__4122\,
            I => \prescale_cntZ0Z_2\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4119\,
            I => \prescale_cntZ0Z_2\
        );

    \I__815\ : InMux
    port map (
            O => \N__4114\,
            I => \N__4111\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4111\,
            I => \prescale_cnt_p1Z0Z_2\
        );

    \I__813\ : InMux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__811\ : Span4Mux_h
    port map (
            O => \N__4102\,
            I => \N__4098\
        );

    \I__810\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4095\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__4098\,
            I => \prescale_cntZ0Z_13\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4095\,
            I => \prescale_cntZ0Z_13\
        );

    \I__807\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4087\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_1\
        );

    \I__805\ : InMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__4075\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_11\
        );

    \I__801\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4069\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_16\
        );

    \I__799\ : InMux
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__797\ : Span4Mux_v
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__4057\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_21\
        );

    \I__795\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4051\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__4051\,
            I => \N__4048\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__4048\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_31\
        );

    \I__792\ : InMux
    port map (
            O => \N__4045\,
            I => proc_pwm_cnt_prescale_cnt10
        );

    \I__791\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4036\
        );

    \I__790\ : InMux
    port map (
            O => \N__4041\,
            I => \N__4036\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4036\,
            I => \N__4033\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4033\,
            I => \proc_pwm_cnt_prescale_cnt10_THRU_CO\
        );

    \I__787\ : InMux
    port map (
            O => \N__4030\,
            I => \N__4027\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4027\,
            I => \N__4024\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__4024\,
            I => pwm_prescale_c_1
        );

    \I__784\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4018\,
            I => \N__4015\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__4015\,
            I => \N__4012\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__4012\,
            I => \N__4009\
        );

    \I__780\ : Sp12to4
    port map (
            O => \N__4009\,
            I => \N__4006\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__4006\,
            I => pwm_lout_c_5
        );

    \I__778\ : InMux
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4000\,
            I => \N__3997\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__3997\,
            I => \pwm_lout_p1Z0Z_5\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__774\ : InMux
    port map (
            O => \N__3991\,
            I => \N__3988\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3988\,
            I => \prescale_stop_p1Z0Z_8\
        );

    \I__772\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__3979\,
            I => \N__3975\
        );

    \I__769\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__3975\,
            I => \prescale_cntZ0Z_8\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__3972\,
            I => \prescale_cntZ0Z_8\
        );

    \I__766\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3964\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__3964\,
            I => \prescale_cnt_p1Z0Z_8\
        );

    \I__764\ : InMux
    port map (
            O => \N__3961\,
            I => \N__3958\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__3958\,
            I => \N__3955\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__3955\,
            I => \N__3951\
        );

    \I__761\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3948\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3951\,
            I => \prescale_cntZ0Z_9\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3948\,
            I => \prescale_cntZ0Z_9\
        );

    \I__758\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3940\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__3940\,
            I => \prescale_cnt_p1Z0Z_9\
        );

    \I__756\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3931\
        );

    \I__755\ : InMux
    port map (
            O => \N__3936\,
            I => \N__3931\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__3931\,
            I => \prescale_stop_p1Z0Z_2\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__3928\,
            I => \N__3925\
        );

    \I__752\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3922\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__3922\,
            I => \prescale_stop_p1Z0Z_3\
        );

    \I__750\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3916\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__3916\,
            I => \N__3913\
        );

    \I__748\ : Span4Mux_h
    port map (
            O => \N__3913\,
            I => \N__3910\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__3910\,
            I => \proc_pwm_cnt_prescale_cnt10_0_N_41\
        );

    \I__746\ : CascadeMux
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__745\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__3901\,
            I => \prescale_stop_p1Z0Z_1\
        );

    \I__743\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3895\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__3895\,
            I => \N__3892\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__3892\,
            I => \N__3889\
        );

    \I__740\ : Span4Mux_v
    port map (
            O => \N__3889\,
            I => \N__3886\
        );

    \I__739\ : Span4Mux_v
    port map (
            O => \N__3886\,
            I => \N__3883\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__3883\,
            I => pwm_lout_c_4
        );

    \I__737\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3877\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3877\,
            I => \N__3874\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__3874\,
            I => \pwm_lout_p1Z0Z_4\
        );

    \I__734\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3868\,
            I => \N__3865\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__3865\,
            I => \N__3861\
        );

    \I__731\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3858\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__3861\,
            I => \prescale_cntZ0Z_5\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__3858\,
            I => \prescale_cntZ0Z_5\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__3853\,
            I => \N__3850\
        );

    \I__727\ : InMux
    port map (
            O => \N__3850\,
            I => \N__3847\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__3847\,
            I => \prescale_stop_p1Z0Z_15\
        );

    \I__725\ : InMux
    port map (
            O => \N__3844\,
            I => \N__3841\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__723\ : Span12Mux_v
    port map (
            O => \N__3838\,
            I => \N__3834\
        );

    \I__722\ : InMux
    port map (
            O => \N__3837\,
            I => \N__3831\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__3834\,
            I => \prescale_cntZ0Z_14\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3831\,
            I => \prescale_cntZ0Z_14\
        );

    \I__719\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3823\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__3823\,
            I => \prescale_cnt_p1Z0Z_14\
        );

    \I__717\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3817\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3817\,
            I => \N__3814\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__3814\,
            I => \N__3811\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__3811\,
            I => \N__3807\
        );

    \I__713\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3804\
        );

    \I__712\ : Odrv4
    port map (
            O => \N__3807\,
            I => \prescale_cntZ0Z_15\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__3804\,
            I => \prescale_cntZ0Z_15\
        );

    \I__710\ : InMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3796\,
            I => \prescale_cnt_p1Z0Z_15\
        );

    \I__708\ : InMux
    port map (
            O => \N__3793\,
            I => prescale_cnt_cry_8
        );

    \I__707\ : InMux
    port map (
            O => \N__3790\,
            I => \N__3787\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3787\,
            I => \N__3783\
        );

    \I__705\ : InMux
    port map (
            O => \N__3786\,
            I => \N__3780\
        );

    \I__704\ : Odrv12
    port map (
            O => \N__3783\,
            I => \prescale_cntZ0Z_10\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3780\,
            I => \prescale_cntZ0Z_10\
        );

    \I__702\ : InMux
    port map (
            O => \N__3775\,
            I => prescale_cnt_cry_9
        );

    \I__701\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3769\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3769\,
            I => \N__3765\
        );

    \I__699\ : InMux
    port map (
            O => \N__3768\,
            I => \N__3762\
        );

    \I__698\ : Odrv12
    port map (
            O => \N__3765\,
            I => \prescale_cntZ0Z_11\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3762\,
            I => \prescale_cntZ0Z_11\
        );

    \I__696\ : InMux
    port map (
            O => \N__3757\,
            I => prescale_cnt_cry_10
        );

    \I__695\ : InMux
    port map (
            O => \N__3754\,
            I => prescale_cnt_cry_11
        );

    \I__694\ : InMux
    port map (
            O => \N__3751\,
            I => prescale_cnt_cry_12
        );

    \I__693\ : InMux
    port map (
            O => \N__3748\,
            I => prescale_cnt_cry_13
        );

    \I__692\ : InMux
    port map (
            O => \N__3745\,
            I => prescale_cnt_cry_14
        );

    \I__691\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3724\
        );

    \I__690\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3715\
        );

    \I__689\ : InMux
    port map (
            O => \N__3740\,
            I => \N__3715\
        );

    \I__688\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3715\
        );

    \I__687\ : InMux
    port map (
            O => \N__3738\,
            I => \N__3715\
        );

    \I__686\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3706\
        );

    \I__685\ : InMux
    port map (
            O => \N__3736\,
            I => \N__3706\
        );

    \I__684\ : InMux
    port map (
            O => \N__3735\,
            I => \N__3706\
        );

    \I__683\ : InMux
    port map (
            O => \N__3734\,
            I => \N__3706\
        );

    \I__682\ : InMux
    port map (
            O => \N__3733\,
            I => \N__3699\
        );

    \I__681\ : InMux
    port map (
            O => \N__3732\,
            I => \N__3699\
        );

    \I__680\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3699\
        );

    \I__679\ : InMux
    port map (
            O => \N__3730\,
            I => \N__3690\
        );

    \I__678\ : InMux
    port map (
            O => \N__3729\,
            I => \N__3690\
        );

    \I__677\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3690\
        );

    \I__676\ : InMux
    port map (
            O => \N__3727\,
            I => \N__3690\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__3724\,
            I => \N_8\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3715\,
            I => \N_8\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__3706\,
            I => \N_8\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3699\,
            I => \N_8\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N_8\
        );

    \I__670\ : InMux
    port map (
            O => \N__3679\,
            I => \bfn_3_14_0_\
        );

    \I__669\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3668\
        );

    \I__668\ : InMux
    port map (
            O => \N__3675\,
            I => \N__3668\
        );

    \I__667\ : InMux
    port map (
            O => \N__3674\,
            I => \N__3663\
        );

    \I__666\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3663\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3668\,
            I => \prescale_stop_p1Z0Z_0\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3663\,
            I => \prescale_stop_p1Z0Z_0\
        );

    \I__663\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3654\
        );

    \I__662\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3651\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3654\,
            I => \prescale_cntZ0Z_1\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3651\,
            I => \prescale_cntZ0Z_1\
        );

    \I__659\ : InMux
    port map (
            O => \N__3646\,
            I => prescale_cnt_cry_0
        );

    \I__658\ : InMux
    port map (
            O => \N__3643\,
            I => prescale_cnt_cry_1
        );

    \I__657\ : InMux
    port map (
            O => \N__3640\,
            I => prescale_cnt_cry_2
        );

    \I__656\ : InMux
    port map (
            O => \N__3637\,
            I => prescale_cnt_cry_3
        );

    \I__655\ : InMux
    port map (
            O => \N__3634\,
            I => prescale_cnt_cry_4
        );

    \I__654\ : InMux
    port map (
            O => \N__3631\,
            I => \N__3628\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3628\,
            I => \N__3624\
        );

    \I__652\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__3624\,
            I => \prescale_cntZ0Z_6\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__3621\,
            I => \prescale_cntZ0Z_6\
        );

    \I__649\ : InMux
    port map (
            O => \N__3616\,
            I => prescale_cnt_cry_5
        );

    \I__648\ : InMux
    port map (
            O => \N__3613\,
            I => \N__3610\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3610\,
            I => \N__3606\
        );

    \I__646\ : InMux
    port map (
            O => \N__3609\,
            I => \N__3603\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__3606\,
            I => \prescale_cntZ0Z_7\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3603\,
            I => \prescale_cntZ0Z_7\
        );

    \I__643\ : InMux
    port map (
            O => \N__3598\,
            I => prescale_cnt_cry_6
        );

    \I__642\ : InMux
    port map (
            O => \N__3595\,
            I => \bfn_3_13_0_\
        );

    \I__641\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3588\
        );

    \I__640\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3585\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__3588\,
            I => \N__3580\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3580\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__3580\,
            I => \pwm_ctrl_p1Z0Z_0\
        );

    \I__636\ : InMux
    port map (
            O => \N__3577\,
            I => \N__3573\
        );

    \I__635\ : InMux
    port map (
            O => \N__3576\,
            I => \N__3570\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3573\,
            I => \N__3567\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3570\,
            I => \N__3564\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3567\,
            I => \pwm_ctrl_p1Z0Z_1\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3564\,
            I => \pwm_ctrl_p1Z0Z_1\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__3559\,
            I => \pwm_loc_1_sqmuxa_cascade_\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3556\,
            I => \un1_pwm_loc8_1_0_cascade_\
        );

    \I__628\ : CEMux
    port map (
            O => \N__3553\,
            I => \N__3549\
        );

    \I__627\ : CEMux
    port map (
            O => \N__3552\,
            I => \N__3546\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__3549\,
            I => pwm_cnte_0_i
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3546\,
            I => pwm_cnte_0_i
        );

    \I__624\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3538\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3538\,
            I => un1_pwm_loc8_1_0
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3535\,
            I => \N__3531\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__3534\,
            I => \N__3526\
        );

    \I__620\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3519\
        );

    \I__619\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3519\
        );

    \I__618\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3519\
        );

    \I__617\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3516\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3519\,
            I => \N__3513\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3516\,
            I => \N__3510\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__3513\,
            I => \prescale_tickZ0\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3510\,
            I => \prescale_tickZ0\
        );

    \I__612\ : InMux
    port map (
            O => \N__3505\,
            I => \N__3502\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__3502\,
            I => pwm_loc_1_sqmuxa
        );

    \I__610\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3496\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3496\,
            I => pwm_loc_0_sqmuxa_1
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__3493\,
            I => \pwm_loc_1_sqmuxa_1_cascade_\
        );

    \I__607\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3487\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__605\ : Span4Mux_h
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__3481\,
            I => \N__3477\
        );

    \I__603\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3474\
        );

    \I__602\ : Odrv4
    port map (
            O => \N__3477\,
            I => \pwm_locZ0\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__3474\,
            I => \pwm_locZ0\
        );

    \I__600\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3464\
        );

    \I__599\ : InMux
    port map (
            O => \N__3468\,
            I => \N__3459\
        );

    \I__598\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3459\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3464\,
            I => \proc_pwm_fsm_pwm_loc20_THRU_CO\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3459\,
            I => \proc_pwm_fsm_pwm_loc20_THRU_CO\
        );

    \I__595\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3451\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__3451\,
            I => \N_87\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__3448\,
            I => \N__3445\
        );

    \I__592\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3437\
        );

    \I__591\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3434\
        );

    \I__590\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3425\
        );

    \I__589\ : InMux
    port map (
            O => \N__3442\,
            I => \N__3425\
        );

    \I__588\ : InMux
    port map (
            O => \N__3441\,
            I => \N__3425\
        );

    \I__587\ : InMux
    port map (
            O => \N__3440\,
            I => \N__3425\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__3437\,
            I => \pwm_toglZ0\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3434\,
            I => \pwm_toglZ0\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3425\,
            I => \pwm_toglZ0\
        );

    \I__583\ : InMux
    port map (
            O => \N__3418\,
            I => \N__3406\
        );

    \I__582\ : InMux
    port map (
            O => \N__3417\,
            I => \N__3406\
        );

    \I__581\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3406\
        );

    \I__580\ : InMux
    port map (
            O => \N__3415\,
            I => \N__3406\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__3406\,
            I => \N__3403\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__3403\,
            I => \N_86\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__3400\,
            I => \N_87_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__3397\,
            I => \N__3388\
        );

    \I__575\ : InMux
    port map (
            O => \N__3396\,
            I => \N__3388\
        );

    \I__574\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3388\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3388\,
            I => \N__3384\
        );

    \I__572\ : InMux
    port map (
            O => \N__3387\,
            I => \N__3381\
        );

    \I__571\ : Span4Mux_h
    port map (
            O => \N__3384\,
            I => \N__3378\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3381\,
            I => \proc_pwm_fsm_pwm_loc8_THRU_CO\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__3378\,
            I => \proc_pwm_fsm_pwm_loc8_THRU_CO\
        );

    \I__568\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3359\
        );

    \I__567\ : InMux
    port map (
            O => \N__3372\,
            I => \N__3359\
        );

    \I__566\ : InMux
    port map (
            O => \N__3371\,
            I => \N__3359\
        );

    \I__565\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3359\
        );

    \I__564\ : InMux
    port map (
            O => \N__3369\,
            I => \N__3348\
        );

    \I__563\ : InMux
    port map (
            O => \N__3368\,
            I => \N__3348\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3359\,
            I => \N__3345\
        );

    \I__561\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3340\
        );

    \I__560\ : InMux
    port map (
            O => \N__3357\,
            I => \N__3340\
        );

    \I__559\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3331\
        );

    \I__558\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3331\
        );

    \I__557\ : InMux
    port map (
            O => \N__3354\,
            I => \N__3331\
        );

    \I__556\ : InMux
    port map (
            O => \N__3353\,
            I => \N__3331\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__3348\,
            I => \N_78_0_i\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__3345\,
            I => \N_78_0_i\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3340\,
            I => \N_78_0_i\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3331\,
            I => \N_78_0_i\
        );

    \I__551\ : InMux
    port map (
            O => \N__3322\,
            I => \N__3318\
        );

    \I__550\ : InMux
    port map (
            O => \N__3321\,
            I => \N__3315\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3318\,
            I => \prescale_cntZ0Z_0\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3315\,
            I => \prescale_cntZ0Z_0\
        );

    \I__547\ : InMux
    port map (
            O => \N__3310\,
            I => \N__3307\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3307\,
            I => prescale_cnt_s_0
        );

    \I__545\ : InMux
    port map (
            O => \N__3304\,
            I => \bfn_3_12_0_\
        );

    \I__544\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3298\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3298\,
            I => \prescale_stop_p1Z0Z_6\
        );

    \I__542\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3292\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3292\,
            I => \prescale_cnt_p1Z0Z_7\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__3289\,
            I => \N__3286\
        );

    \I__539\ : InMux
    port map (
            O => \N__3286\,
            I => \N__3283\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3283\,
            I => \prescale_stop_p1Z0Z_7\
        );

    \I__537\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3277\,
            I => \prescale_cnt_p1Z0Z_6\
        );

    \I__535\ : InMux
    port map (
            O => \N__3274\,
            I => \N__3271\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3271\,
            I => \prescale_stop_p1Z0Z_10\
        );

    \I__533\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3265\,
            I => \prescale_cnt_p1Z0Z_11\
        );

    \I__531\ : InMux
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3259\,
            I => \prescale_cnt_p1Z0Z_10\
        );

    \I__529\ : InMux
    port map (
            O => \N__3256\,
            I => \N__3251\
        );

    \I__528\ : InMux
    port map (
            O => \N__3255\,
            I => \N__3248\
        );

    \I__527\ : InMux
    port map (
            O => \N__3254\,
            I => \N__3245\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3251\,
            I => \pwm_cntZ0Z_1\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3248\,
            I => \pwm_cntZ0Z_1\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3245\,
            I => \pwm_cntZ0Z_1\
        );

    \I__523\ : InMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__521\ : Odrv4
    port map (
            O => \N__3232\,
            I => \pwm_lout_p1Z0Z_1\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__3229\,
            I => \N__3225\
        );

    \I__519\ : InMux
    port map (
            O => \N__3228\,
            I => \N__3221\
        );

    \I__518\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3218\
        );

    \I__517\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3215\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3221\,
            I => \pwm_cntZ0Z_0\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3218\,
            I => \pwm_cntZ0Z_0\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3215\,
            I => \pwm_cntZ0Z_0\
        );

    \I__513\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3205\,
            I => \pwm_lout_p1Z0Z_0\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__510\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3196\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3196\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_26\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__3193\,
            I => \N__3189\
        );

    \I__507\ : InMux
    port map (
            O => \N__3192\,
            I => \N__3185\
        );

    \I__506\ : InMux
    port map (
            O => \N__3189\,
            I => \N__3182\
        );

    \I__505\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3179\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3185\,
            I => \pwm_cntZ0Z_5\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3182\,
            I => \pwm_cntZ0Z_5\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3179\,
            I => \pwm_cntZ0Z_5\
        );

    \I__501\ : InMux
    port map (
            O => \N__3172\,
            I => \N__3167\
        );

    \I__500\ : InMux
    port map (
            O => \N__3171\,
            I => \N__3164\
        );

    \I__499\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3161\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3167\,
            I => \pwm_cntZ0Z_4\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3164\,
            I => \pwm_cntZ0Z_4\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3161\,
            I => \pwm_cntZ0Z_4\
        );

    \I__495\ : CascadeMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__494\ : InMux
    port map (
            O => \N__3151\,
            I => \N__3148\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3148\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_16\
        );

    \I__492\ : InMux
    port map (
            O => \N__3145\,
            I => \N__3142\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__490\ : Span4Mux_h
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__3130\,
            I => pwm_lout_c_11
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__485\ : InMux
    port map (
            O => \N__3124\,
            I => \N__3121\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3121\,
            I => \pwm_lout_p1Z0Z_11\
        );

    \I__483\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3115\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3115\,
            I => \N__3112\
        );

    \I__481\ : Span12Mux_v
    port map (
            O => \N__3112\,
            I => \N__3109\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__3109\,
            I => pwm_lout_c_10
        );

    \I__479\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3103\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3103\,
            I => \pwm_lout_p1Z0Z_10\
        );

    \I__477\ : InMux
    port map (
            O => \N__3100\,
            I => \N__3097\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3097\,
            I => \N__3094\
        );

    \I__475\ : Sp12to4
    port map (
            O => \N__3094\,
            I => \N__3091\
        );

    \I__474\ : Span12Mux_v
    port map (
            O => \N__3091\,
            I => \N__3088\
        );

    \I__473\ : Odrv12
    port map (
            O => \N__3088\,
            I => pwm_lout_c_1
        );

    \I__472\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3082\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__470\ : Span4Mux_v
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__469\ : Sp12to4
    port map (
            O => \N__3076\,
            I => \N__3073\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__3073\,
            I => pwm_ctrl_c_1
        );

    \I__467\ : InMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3064\
        );

    \I__465\ : Span12Mux_h
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__464\ : Span12Mux_v
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__463\ : Odrv12
    port map (
            O => \N__3058\,
            I => pwm_lout_c_0
        );

    \I__462\ : InMux
    port map (
            O => \N__3055\,
            I => pwm_cnt_cry_9
        );

    \I__461\ : InMux
    port map (
            O => \N__3052\,
            I => pwm_cnt_cry_10
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3049\,
            I => \N_8_cascade_\
        );

    \I__459\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3043\,
            I => \prescale_cnt_p1Z0Z_0\
        );

    \I__457\ : InMux
    port map (
            O => \N__3040\,
            I => \N__3037\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3037\,
            I => \prescale_cnt_p1Z0Z_1\
        );

    \I__455\ : InMux
    port map (
            O => \N__3034\,
            I => \N__3025\
        );

    \I__454\ : InMux
    port map (
            O => \N__3033\,
            I => \N__3025\
        );

    \I__453\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3025\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3025\,
            I => \N_38\
        );

    \I__451\ : InMux
    port map (
            O => \N__3022\,
            I => \N__3017\
        );

    \I__450\ : InMux
    port map (
            O => \N__3021\,
            I => \N__3014\
        );

    \I__449\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3011\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3017\,
            I => \N__3008\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3014\,
            I => \pwm_cntZ0Z_11\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3011\,
            I => \pwm_cntZ0Z_11\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__3008\,
            I => \pwm_cntZ0Z_11\
        );

    \I__444\ : InMux
    port map (
            O => \N__3001\,
            I => \N__2996\
        );

    \I__443\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2993\
        );

    \I__442\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2990\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__2996\,
            I => \N__2987\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__2993\,
            I => \pwm_cntZ0Z_10\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__2990\,
            I => \pwm_cntZ0Z_10\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__2987\,
            I => \pwm_cntZ0Z_10\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__2980\,
            I => \N__2977\
        );

    \I__436\ : InMux
    port map (
            O => \N__2977\,
            I => \N__2974\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2974\,
            I => \N__2971\
        );

    \I__434\ : Odrv12
    port map (
            O => \N__2971\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_1\
        );

    \I__433\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2963\
        );

    \I__432\ : InMux
    port map (
            O => \N__2967\,
            I => \N__2960\
        );

    \I__431\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2957\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__2963\,
            I => \pwm_cntZ0Z_2\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2960\,
            I => \pwm_cntZ0Z_2\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2957\,
            I => \pwm_cntZ0Z_2\
        );

    \I__427\ : InMux
    port map (
            O => \N__2950\,
            I => pwm_cnt_cry_1
        );

    \I__426\ : InMux
    port map (
            O => \N__2947\,
            I => \N__2942\
        );

    \I__425\ : InMux
    port map (
            O => \N__2946\,
            I => \N__2937\
        );

    \I__424\ : InMux
    port map (
            O => \N__2945\,
            I => \N__2937\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__2942\,
            I => \pwm_cntZ0Z_3\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2937\,
            I => \pwm_cntZ0Z_3\
        );

    \I__421\ : InMux
    port map (
            O => \N__2932\,
            I => pwm_cnt_cry_2
        );

    \I__420\ : InMux
    port map (
            O => \N__2929\,
            I => pwm_cnt_cry_3
        );

    \I__419\ : InMux
    port map (
            O => \N__2926\,
            I => pwm_cnt_cry_4
        );

    \I__418\ : InMux
    port map (
            O => \N__2923\,
            I => \N__2918\
        );

    \I__417\ : InMux
    port map (
            O => \N__2922\,
            I => \N__2915\
        );

    \I__416\ : InMux
    port map (
            O => \N__2921\,
            I => \N__2912\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2918\,
            I => \pwm_cntZ0Z_6\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2915\,
            I => \pwm_cntZ0Z_6\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2912\,
            I => \pwm_cntZ0Z_6\
        );

    \I__412\ : InMux
    port map (
            O => \N__2905\,
            I => pwm_cnt_cry_5
        );

    \I__411\ : InMux
    port map (
            O => \N__2902\,
            I => \N__2897\
        );

    \I__410\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2894\
        );

    \I__409\ : InMux
    port map (
            O => \N__2900\,
            I => \N__2891\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2897\,
            I => \pwm_cntZ0Z_7\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2894\,
            I => \pwm_cntZ0Z_7\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2891\,
            I => \pwm_cntZ0Z_7\
        );

    \I__405\ : InMux
    port map (
            O => \N__2884\,
            I => pwm_cnt_cry_6
        );

    \I__404\ : InMux
    port map (
            O => \N__2881\,
            I => \N__2876\
        );

    \I__403\ : InMux
    port map (
            O => \N__2880\,
            I => \N__2873\
        );

    \I__402\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2870\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2876\,
            I => \N__2867\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2873\,
            I => \pwm_cntZ0Z_8\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2870\,
            I => \pwm_cntZ0Z_8\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__2867\,
            I => \pwm_cntZ0Z_8\
        );

    \I__397\ : InMux
    port map (
            O => \N__2860\,
            I => \bfn_2_12_0_\
        );

    \I__396\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2852\
        );

    \I__395\ : InMux
    port map (
            O => \N__2856\,
            I => \N__2849\
        );

    \I__394\ : InMux
    port map (
            O => \N__2855\,
            I => \N__2846\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2852\,
            I => \N__2843\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2849\,
            I => \pwm_cntZ0Z_9\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2846\,
            I => \pwm_cntZ0Z_9\
        );

    \I__390\ : Odrv4
    port map (
            O => \N__2843\,
            I => \pwm_cntZ0Z_9\
        );

    \I__389\ : InMux
    port map (
            O => \N__2836\,
            I => pwm_cnt_cry_8
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2833\,
            I => \N__2830\
        );

    \I__387\ : InMux
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2827\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_21\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__2824\,
            I => \N__2821\
        );

    \I__384\ : InMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2818\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_6\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2815\,
            I => \N__2812\
        );

    \I__381\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2809\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2809\,
            I => \proc_pwm_fsm_pwm_loc20_0_N_11\
        );

    \I__379\ : InMux
    port map (
            O => \N__2806\,
            I => proc_pwm_fsm_pwm_loc20
        );

    \I__378\ : InMux
    port map (
            O => \N__2803\,
            I => \bfn_2_11_0_\
        );

    \I__377\ : InMux
    port map (
            O => \N__2800\,
            I => pwm_cnt_cry_0
        );

    \I__376\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2794\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__2794\,
            I => \N__2791\
        );

    \I__374\ : Span4Mux_v
    port map (
            O => \N__2791\,
            I => \N__2788\
        );

    \I__373\ : Span4Mux_v
    port map (
            O => \N__2788\,
            I => \N__2785\
        );

    \I__372\ : Span4Mux_h
    port map (
            O => \N__2785\,
            I => \N__2782\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__2782\,
            I => pwm_hout_c_7
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__369\ : InMux
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__367\ : Span4Mux_h
    port map (
            O => \N__2770\,
            I => \N__2767\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__2767\,
            I => \pwm_hout_p1Z0Z_7\
        );

    \I__365\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2761\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__363\ : Span4Mux_h
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__362\ : Span4Mux_v
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__2749\,
            I => pwm_hout_c_11
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__2746\,
            I => \N__2743\
        );

    \I__358\ : InMux
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__357\ : LocalMux
    port map (
            O => \N__2740\,
            I => \pwm_hout_p1Z0Z_11\
        );

    \I__356\ : InMux
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__354\ : Span4Mux_v
    port map (
            O => \N__2731\,
            I => \N__2728\
        );

    \I__353\ : Span4Mux_h
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__352\ : Odrv4
    port map (
            O => \N__2725\,
            I => pwm_prescale_c_0
        );

    \I__351\ : InMux
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2719\,
            I => \N__2716\
        );

    \I__349\ : Span4Mux_v
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__348\ : Sp12to4
    port map (
            O => \N__2713\,
            I => \N__2710\
        );

    \I__347\ : Odrv12
    port map (
            O => \N__2710\,
            I => pwm_lout_c_7
        );

    \I__346\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2704\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__2704\,
            I => \N__2701\
        );

    \I__344\ : Odrv12
    port map (
            O => \N__2701\,
            I => \pwm_lout_p1Z0Z_7\
        );

    \I__343\ : InMux
    port map (
            O => \N__2698\,
            I => \N__2695\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__2695\,
            I => \N__2692\
        );

    \I__341\ : Span12Mux_v
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__340\ : Odrv12
    port map (
            O => \N__2689\,
            I => pwm_prescale_c_2
        );

    \I__339\ : InMux
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2683\,
            I => \N__2680\
        );

    \I__337\ : Span12Mux_v
    port map (
            O => \N__2680\,
            I => \N__2677\
        );

    \I__336\ : Odrv12
    port map (
            O => \N__2677\,
            I => pwm_lout_c_8
        );

    \I__335\ : InMux
    port map (
            O => \N__2674\,
            I => \N__2671\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2671\,
            I => \N__2668\
        );

    \I__333\ : Span12Mux_v
    port map (
            O => \N__2668\,
            I => \N__2665\
        );

    \I__332\ : Odrv12
    port map (
            O => \N__2665\,
            I => pwm_ctrl_c_0
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__330\ : InMux
    port map (
            O => \N__2659\,
            I => \N__2656\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2656\,
            I => \pwm_lout_p1Z0Z_8\
        );

    \I__328\ : InMux
    port map (
            O => \N__2653\,
            I => \N__2650\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__2650\,
            I => \pwm_lout_p1Z0Z_9\
        );

    \I__326\ : InMux
    port map (
            O => \N__2647\,
            I => \N__2644\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__2644\,
            I => \N__2641\
        );

    \I__324\ : Span4Mux_h
    port map (
            O => \N__2641\,
            I => \N__2638\
        );

    \I__323\ : Span4Mux_v
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__322\ : Odrv4
    port map (
            O => \N__2635\,
            I => pwm_hout_c_0
        );

    \I__321\ : InMux
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2629\,
            I => \pwm_hout_p1Z0Z_0\
        );

    \I__319\ : InMux
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2623\,
            I => \N__2620\
        );

    \I__317\ : Span4Mux_v
    port map (
            O => \N__2620\,
            I => \N__2617\
        );

    \I__316\ : Span4Mux_h
    port map (
            O => \N__2617\,
            I => \N__2614\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__2614\,
            I => pwm_hout_c_3
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2611\,
            I => \N__2608\
        );

    \I__313\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2605\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__2605\,
            I => \pwm_hout_p1Z0Z_3\
        );

    \I__311\ : InMux
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__309\ : Span12Mux_h
    port map (
            O => \N__2596\,
            I => \N__2593\
        );

    \I__308\ : Span12Mux_v
    port map (
            O => \N__2593\,
            I => \N__2590\
        );

    \I__307\ : Odrv12
    port map (
            O => \N__2590\,
            I => pwm_lout_c_2
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__305\ : InMux
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2581\,
            I => \pwm_lout_p1Z0Z_2\
        );

    \I__303\ : InMux
    port map (
            O => \N__2578\,
            I => \N__2575\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2575\,
            I => \N__2572\
        );

    \I__301\ : Span4Mux_h
    port map (
            O => \N__2572\,
            I => \N__2569\
        );

    \I__300\ : Span4Mux_v
    port map (
            O => \N__2569\,
            I => \N__2566\
        );

    \I__299\ : Odrv4
    port map (
            O => \N__2566\,
            I => pwm_hout_c_1
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__2563\,
            I => \N__2560\
        );

    \I__297\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2557\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2557\,
            I => \pwm_hout_p1Z0Z_1\
        );

    \I__295\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2551\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2551\,
            I => \N__2548\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__2548\,
            I => \N__2545\
        );

    \I__292\ : Span4Mux_v
    port map (
            O => \N__2545\,
            I => \N__2542\
        );

    \I__291\ : Span4Mux_h
    port map (
            O => \N__2542\,
            I => \N__2539\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__2539\,
            I => pwm_hout_c_2
        );

    \I__289\ : InMux
    port map (
            O => \N__2536\,
            I => \N__2533\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2533\,
            I => \pwm_hout_p1Z0Z_2\
        );

    \I__287\ : InMux
    port map (
            O => \N__2530\,
            I => \N__2527\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__2527\,
            I => \N__2524\
        );

    \I__285\ : Odrv12
    port map (
            O => \N__2524\,
            I => pwm_lout_c_3
        );

    \I__284\ : InMux
    port map (
            O => \N__2521\,
            I => \N__2518\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2518\,
            I => \pwm_lout_p1Z0Z_3\
        );

    \I__282\ : InMux
    port map (
            O => \N__2515\,
            I => \N__2512\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2512\,
            I => \N__2509\
        );

    \I__280\ : Odrv12
    port map (
            O => \N__2509\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_1\
        );

    \I__279\ : InMux
    port map (
            O => \N__2506\,
            I => \N__2503\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2503\,
            I => \N__2500\
        );

    \I__277\ : Sp12to4
    port map (
            O => \N__2500\,
            I => \N__2497\
        );

    \I__276\ : Span12Mux_v
    port map (
            O => \N__2497\,
            I => \N__2494\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__2494\,
            I => pwm_hout_c_6
        );

    \I__274\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2488\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2488\,
            I => \N__2485\
        );

    \I__272\ : Odrv4
    port map (
            O => \N__2485\,
            I => \pwm_hout_p1Z0Z_6\
        );

    \I__271\ : InMux
    port map (
            O => \N__2482\,
            I => \N__2479\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2479\,
            I => \N__2476\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__2476\,
            I => \N__2473\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__2473\,
            I => \N__2470\
        );

    \I__267\ : Span4Mux_h
    port map (
            O => \N__2470\,
            I => \N__2467\
        );

    \I__266\ : Odrv4
    port map (
            O => \N__2467\,
            I => pwm_hout_c_10
        );

    \I__265\ : InMux
    port map (
            O => \N__2464\,
            I => \N__2461\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2461\,
            I => \pwm_hout_p1Z0Z_10\
        );

    \I__263\ : CascadeMux
    port map (
            O => \N__2458\,
            I => \N__2455\
        );

    \I__262\ : InMux
    port map (
            O => \N__2455\,
            I => \N__2452\
        );

    \I__261\ : LocalMux
    port map (
            O => \N__2452\,
            I => \pwm_lout_p1Z0Z_6\
        );

    \I__260\ : CascadeMux
    port map (
            O => \N__2449\,
            I => \N__2446\
        );

    \I__259\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2443\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__2443\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_26\
        );

    \I__257\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2437\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2437\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_6\
        );

    \I__255\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2431\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__2431\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_16\
        );

    \I__253\ : InMux
    port map (
            O => \N__2428\,
            I => \N__2425\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2425\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_21\
        );

    \I__251\ : InMux
    port map (
            O => \N__2422\,
            I => \N__2419\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2419\,
            I => \N__2416\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__2416\,
            I => \pwm_hout_p1Z0Z_8\
        );

    \I__248\ : CascadeMux
    port map (
            O => \N__2413\,
            I => \N__2410\
        );

    \I__247\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2407\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__2407\,
            I => \N__2404\
        );

    \I__245\ : Span4Mux_v
    port map (
            O => \N__2404\,
            I => \N__2401\
        );

    \I__244\ : Odrv4
    port map (
            O => \N__2401\,
            I => \pwm_hout_p1Z0Z_9\
        );

    \I__243\ : InMux
    port map (
            O => \N__2398\,
            I => \N__2395\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2395\,
            I => \proc_pwm_fsm_pwm_loc8_0_N_11\
        );

    \I__241\ : InMux
    port map (
            O => \N__2392\,
            I => \N__2389\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2389\,
            I => \N__2386\
        );

    \I__239\ : Span4Mux_v
    port map (
            O => \N__2386\,
            I => \N__2383\
        );

    \I__238\ : Sp12to4
    port map (
            O => \N__2383\,
            I => \N__2380\
        );

    \I__237\ : Span12Mux_h
    port map (
            O => \N__2380\,
            I => \N__2377\
        );

    \I__236\ : Odrv12
    port map (
            O => \N__2377\,
            I => pwm_hout_c_5
        );

    \I__235\ : CascadeMux
    port map (
            O => \N__2374\,
            I => \N__2371\
        );

    \I__234\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2368\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2368\,
            I => \pwm_hout_p1Z0Z_5\
        );

    \I__232\ : InMux
    port map (
            O => \N__2365\,
            I => \N__2362\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2362\,
            I => \N__2359\
        );

    \I__230\ : Span4Mux_h
    port map (
            O => \N__2359\,
            I => \N__2356\
        );

    \I__229\ : Span4Mux_v
    port map (
            O => \N__2356\,
            I => \N__2353\
        );

    \I__228\ : Span4Mux_v
    port map (
            O => \N__2353\,
            I => \N__2350\
        );

    \I__227\ : Span4Mux_v
    port map (
            O => \N__2350\,
            I => \N__2347\
        );

    \I__226\ : Odrv4
    port map (
            O => \N__2347\,
            I => pwm_hout_c_4
        );

    \I__225\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2341\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2341\,
            I => \pwm_hout_p1Z0Z_4\
        );

    \I__223\ : InMux
    port map (
            O => \N__2338\,
            I => \N__2335\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2335\,
            I => \N__2332\
        );

    \I__221\ : Sp12to4
    port map (
            O => \N__2332\,
            I => \N__2329\
        );

    \I__220\ : Span12Mux_v
    port map (
            O => \N__2329\,
            I => \N__2326\
        );

    \I__219\ : Odrv12
    port map (
            O => \N__2326\,
            I => pwm_hout_c_9
        );

    \I__218\ : InMux
    port map (
            O => \N__2323\,
            I => \N__2320\
        );

    \I__217\ : LocalMux
    port map (
            O => \N__2320\,
            I => \N__2317\
        );

    \I__216\ : Span4Mux_v
    port map (
            O => \N__2317\,
            I => \N__2314\
        );

    \I__215\ : Span4Mux_v
    port map (
            O => \N__2314\,
            I => \N__2311\
        );

    \I__214\ : Span4Mux_v
    port map (
            O => \N__2311\,
            I => \N__2308\
        );

    \I__213\ : Sp12to4
    port map (
            O => \N__2308\,
            I => \N__2305\
        );

    \I__212\ : Odrv12
    port map (
            O => \N__2305\,
            I => pwm_hout_c_8
        );

    \I__211\ : InMux
    port map (
            O => \N__2302\,
            I => proc_pwm_fsm_pwm_loc8
        );

    \I__210\ : IoInMux
    port map (
            O => \N__2299\,
            I => \N__2296\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__2296\,
            I => \N__2293\
        );

    \I__208\ : IoSpan4Mux
    port map (
            O => \N__2293\,
            I => \N__2290\
        );

    \I__207\ : Span4Mux_s3_h
    port map (
            O => \N__2290\,
            I => \N__2287\
        );

    \I__206\ : Odrv4
    port map (
            O => \N__2287\,
            I => pwm_pin_c
        );

    \I__205\ : InMux
    port map (
            O => \N__2284\,
            I => \N__2281\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__2281\,
            I => \N__2278\
        );

    \I__203\ : Span4Mux_v
    port map (
            O => \N__2278\,
            I => \N__2275\
        );

    \I__202\ : Span4Mux_v
    port map (
            O => \N__2275\,
            I => \N__2272\
        );

    \I__201\ : Sp12to4
    port map (
            O => \N__2272\,
            I => \N__2269\
        );

    \I__200\ : Odrv12
    port map (
            O => \N__2269\,
            I => pwm_lout_c_9
        );

    \I__199\ : InMux
    port map (
            O => \N__2266\,
            I => \N__2263\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__2263\,
            I => \N__2260\
        );

    \I__197\ : Span4Mux_h
    port map (
            O => \N__2260\,
            I => \N__2257\
        );

    \I__196\ : Sp12to4
    port map (
            O => \N__2257\,
            I => \N__2254\
        );

    \I__195\ : Span12Mux_v
    port map (
            O => \N__2254\,
            I => \N__2251\
        );

    \I__194\ : Odrv12
    port map (
            O => \N__2251\,
            I => pwm_lout_c_6
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_7,
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => pwm_cnt_cry_7,
            carryinitout => \bfn_2_12_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => prescale_cnt_cry_7,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_3_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => prescale_cnt_cry_15,
            carryinitout => \bfn_3_14_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \pwm_pinZ0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3490\,
            lcout => pwm_pin_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4393\,
            ce => 'H',
            sr => \N__4317\
        );

    \pwm_lout_p1_9_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2284\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_lout_p1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4385\,
            ce => 'H',
            sr => \N__4308\
        );

    \pwm_lout_p1_6_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_lout_p1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4384\,
            ce => 'H',
            sr => \N__4306\
        );

    \pwm_hout_p1_9_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2338\,
            lcout => \pwm_hout_p1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4384\,
            ce => 'H',
            sr => \N__4306\
        );

    \pwm_hout_p1_8_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2323\,
            lcout => \pwm_hout_p1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4384\,
            ce => 'H',
            sr => \N__4306\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_1_c_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2449\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => proc_pwm_fsm_pwm_loc8_0_data_tmp_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_9_c_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2428\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc8_0_data_tmp_0,
            carryout => proc_pwm_fsm_pwm_loc8_0_data_tmp_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_15_c_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2434\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc8_0_data_tmp_1,
            carryout => proc_pwm_fsm_pwm_loc8_0_data_tmp_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_27_c_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2440\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc8_0_data_tmp_2,
            carryout => proc_pwm_fsm_pwm_loc8_0_data_tmp_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_21_c_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2398\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc8_0_data_tmp_3,
            carryout => proc_pwm_fsm_pwm_loc8_0_data_tmp_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_33_c_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2515\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc8_0_data_tmp_4,
            carryout => proc_pwm_fsm_pwm_loc8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_THRU_LUT4_0_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2302\,
            lcout => \proc_pwm_fsm_pwm_loc8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_27_c_RNO_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__2707\,
            in1 => \N__2901\,
            in2 => \N__2458\,
            in3 => \N__2921\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_1_c_RNO_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2632\,
            in1 => \N__3254\,
            in2 => \N__2563\,
            in3 => \N__3224\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_27_c_RNO_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2491\,
            in1 => \N__2900\,
            in2 => \N__2779\,
            in3 => \N__2922\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_9_c_RNO_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__2967\,
            in1 => \N__2946\,
            in2 => \N__2587\,
            in3 => \N__2521\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_15_c_RNO_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2344\,
            in1 => \N__3188\,
            in2 => \N__2374\,
            in3 => \N__3171\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_9_c_RNO_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2536\,
            in1 => \N__2945\,
            in2 => \N__2611\,
            in3 => \N__2966\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_21_c_RNO_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2422\,
            in1 => \N__2855\,
            in2 => \N__2413\,
            in3 => \N__2879\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_hout_p1_5_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2392\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_hout_p1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_hout_p1_4_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2365\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_hout_p1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_hout_p1_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2647\,
            lcout => \pwm_hout_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_hout_p1_3_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2626\,
            lcout => \pwm_hout_p1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_lout_p1_2_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_lout_p1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_hout_p1_1_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2578\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_hout_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_hout_p1_2_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_hout_p1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \pwm_lout_p1_3_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2530\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_lout_p1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4386\,
            ce => 'H',
            sr => \N__4304\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_33_c_RNO_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2464\,
            in1 => \N__3020\,
            in2 => \N__2746\,
            in3 => \N__2999\,
            lcout => \proc_pwm_fsm_pwm_loc8_0_N_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_hout_p1_6_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2506\,
            lcout => \pwm_hout_p1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_hout_p1_10_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2482\,
            lcout => \pwm_hout_p1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_hout_p1_7_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2797\,
            lcout => \pwm_hout_p1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_hout_p1_11_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2764\,
            lcout => \pwm_hout_p1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_prescale_p1_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2737\,
            lcout => \pwm_prescale_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_lout_p1_7_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2722\,
            lcout => \pwm_lout_p1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4394\,
            ce => 'H',
            sr => \N__4309\
        );

    \pwm_prescale_p1_2_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2698\,
            lcout => \pwm_prescale_p1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4395\,
            ce => 'H',
            sr => \N__4318\
        );

    \pwm_lout_p1_8_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2686\,
            lcout => \pwm_lout_p1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4388\,
            ce => 'H',
            sr => \N__4313\
        );

    \pwm_ctrl_p1_0_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2674\,
            lcout => \pwm_ctrl_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4388\,
            ce => 'H',
            sr => \N__4313\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_21_c_RNO_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__2857\,
            in1 => \N__2881\,
            in2 => \N__2662\,
            in3 => \N__2653\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_1_c_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3202\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => proc_pwm_fsm_pwm_loc20_0_data_tmp_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_9_c_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2833\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc20_0_data_tmp_0,
            carryout => proc_pwm_fsm_pwm_loc20_0_data_tmp_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_15_c_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3154\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc20_0_data_tmp_1,
            carryout => proc_pwm_fsm_pwm_loc20_0_data_tmp_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_27_c_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2824\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc20_0_data_tmp_2,
            carryout => proc_pwm_fsm_pwm_loc20_0_data_tmp_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_21_c_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2815\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc20_0_data_tmp_3,
            carryout => proc_pwm_fsm_pwm_loc20_0_data_tmp_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_33_c_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2980\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_fsm_pwm_loc20_0_data_tmp_4,
            carryout => proc_pwm_fsm_pwm_loc20,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_THRU_LUT4_0_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2806\,
            lcout => \proc_pwm_fsm_pwm_loc20_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_loc_RNO_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011100000"
        )
    port map (
            in0 => \N__3387\,
            in1 => \N__3444\,
            in2 => \N__3534\,
            in3 => \N__3469\,
            lcout => pwm_loc_0_sqmuxa_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_cnt_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__3370\,
            in1 => \N__3228\,
            in2 => \_gnd_net_\,
            in3 => \N__2803\,
            lcout => \pwm_cntZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => pwm_cnt_cry_0,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3353\,
            in1 => \N__3256\,
            in2 => \_gnd_net_\,
            in3 => \N__2800\,
            lcout => \pwm_cntZ0Z_1\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_0,
            carryout => pwm_cnt_cry_1,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3371\,
            in1 => \N__2968\,
            in2 => \_gnd_net_\,
            in3 => \N__2950\,
            lcout => \pwm_cntZ0Z_2\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_1,
            carryout => pwm_cnt_cry_2,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_3_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3354\,
            in1 => \N__2947\,
            in2 => \_gnd_net_\,
            in3 => \N__2932\,
            lcout => \pwm_cntZ0Z_3\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_2,
            carryout => pwm_cnt_cry_3,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_4_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3372\,
            in1 => \N__3172\,
            in2 => \_gnd_net_\,
            in3 => \N__2929\,
            lcout => \pwm_cntZ0Z_4\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_3,
            carryout => pwm_cnt_cry_4,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_5_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3355\,
            in1 => \N__3192\,
            in2 => \_gnd_net_\,
            in3 => \N__2926\,
            lcout => \pwm_cntZ0Z_5\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_4,
            carryout => pwm_cnt_cry_5,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_6_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3373\,
            in1 => \N__2923\,
            in2 => \_gnd_net_\,
            in3 => \N__2905\,
            lcout => \pwm_cntZ0Z_6\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_5,
            carryout => pwm_cnt_cry_6,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_7_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3356\,
            in1 => \N__2902\,
            in2 => \_gnd_net_\,
            in3 => \N__2884\,
            lcout => \pwm_cntZ0Z_7\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_6,
            carryout => pwm_cnt_cry_7,
            clk => \N__4387\,
            ce => \N__3552\,
            sr => \N__4303\
        );

    \pwm_cnt_8_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3369\,
            in1 => \N__2880\,
            in2 => \_gnd_net_\,
            in3 => \N__2860\,
            lcout => \pwm_cntZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_2_12_0_\,
            carryout => pwm_cnt_cry_8,
            clk => \N__4389\,
            ce => \N__3553\,
            sr => \N__4307\
        );

    \pwm_cnt_9_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3357\,
            in1 => \N__2856\,
            in2 => \_gnd_net_\,
            in3 => \N__2836\,
            lcout => \pwm_cntZ0Z_9\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_8,
            carryout => pwm_cnt_cry_9,
            clk => \N__4389\,
            ce => \N__3553\,
            sr => \N__4307\
        );

    \pwm_cnt_10_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3368\,
            in1 => \N__3000\,
            in2 => \_gnd_net_\,
            in3 => \N__3055\,
            lcout => \pwm_cntZ0Z_10\,
            ltout => OPEN,
            carryin => pwm_cnt_cry_9,
            carryout => pwm_cnt_cry_10,
            clk => \N__4389\,
            ce => \N__3553\,
            sr => \N__4307\
        );

    \pwm_cnt_11_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3358\,
            in1 => \N__3021\,
            in2 => \_gnd_net_\,
            in3 => \N__3052\,
            lcout => \pwm_cntZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4389\,
            ce => \N__3553\,
            sr => \N__4307\
        );

    \prescale_tick_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4042\,
            in1 => \N__3033\,
            in2 => \_gnd_net_\,
            in3 => \N__3675\,
            lcout => \prescale_tickZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4396\,
            ce => 'H',
            sr => \N__4310\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNIRR0O1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__3032\,
            in1 => \N__3674\,
            in2 => \_gnd_net_\,
            in3 => \N__4041\,
            lcout => \N_8\,
            ltout => \N_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__3310\,
            in1 => \N__3034\,
            in2 => \N__3049\,
            in3 => \N__3676\,
            lcout => \prescale_cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4396\,
            ce => 'H',
            sr => \N__4310\
        );

    \prescale_cnt_p1_0_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3322\,
            lcout => \prescale_cnt_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4396\,
            ce => 'H',
            sr => \N__4310\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_1_c_RNO_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3673\,
            in1 => \N__3040\,
            in2 => \N__3907\,
            in3 => \N__3046\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_p1_1_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3658\,
            lcout => \prescale_cnt_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4396\,
            ce => 'H',
            sr => \N__4310\
        );

    \pwm_prescale_p1_RNI1QRQ_0_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4648\,
            in1 => \N__4596\,
            in2 => \_gnd_net_\,
            in3 => \N__4434\,
            lcout => \N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_33_c_RNO_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__3022\,
            in1 => \N__3001\,
            in2 => \N__3127\,
            in3 => \N__3106\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_lout_p1_11_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3145\,
            lcout => \pwm_lout_p1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4405\,
            ce => 'H',
            sr => \N__4323\
        );

    \pwm_lout_p1_10_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3118\,
            lcout => \pwm_lout_p1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4405\,
            ce => 'H',
            sr => \N__4323\
        );

    \pwm_lout_p1_1_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3100\,
            lcout => \pwm_lout_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4397\,
            ce => 'H',
            sr => \N__4319\
        );

    \pwm_ctrl_p1_1_LC_3_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_ctrl_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4397\,
            ce => 'H',
            sr => \N__4319\
        );

    \prescale_cnt_p1_11_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3772\,
            lcout => \prescale_cnt_p1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \pwm_lout_p1_0_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_lout_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_cnt_p1_10_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \prescale_cnt_p1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_stop_p1_6_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__4491\,
            in1 => \_gnd_net_\,
            in2 => \N__4603\,
            in3 => \N__4667\,
            lcout => \prescale_stop_p1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_cnt_p1_7_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3613\,
            lcout => \prescale_cnt_p1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_cnt_p1_6_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3631\,
            lcout => \prescale_cnt_p1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_stop_p1_10_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__4666\,
            in1 => \N__4599\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => \prescale_stop_p1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \prescale_stop_p1_7_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4665\,
            lcout => \prescale_stop_p1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4390\,
            ce => 'H',
            sr => \N__4314\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_39_c_RNO_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3301\,
            in1 => \N__3295\,
            in2 => \N__3289\,
            in3 => \N__3280\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_27_c_RNO_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__3274\,
            in1 => \N__3268\,
            in2 => \_gnd_net_\,
            in3 => \N__3262\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_1_c_RNO_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__3255\,
            in1 => \N__3238\,
            in2 => \N__3229\,
            in3 => \N__3208\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctrl_p1_RNI1IE6_0_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3577\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3592\,
            lcout => \N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_15_c_RNO_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__4003\,
            in1 => \N__3880\,
            in2 => \N__3193\,
            in3 => \N__3170\,
            lcout => \proc_pwm_fsm_pwm_loc20_0_N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_ctrl_p1_RNICQ6G_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3591\,
            in1 => \N__3576\,
            in2 => \_gnd_net_\,
            in3 => \N__3467\,
            lcout => pwm_loc_1_sqmuxa,
            ltout => \pwm_loc_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIMT131_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__3441\,
            in1 => \_gnd_net_\,
            in2 => \N__3559\,
            in3 => \N__3395\,
            lcout => un1_pwm_loc8_1_0,
            ltout => \un1_pwm_loc8_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_tick_RNI46OT1_LC_3_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011101110"
        )
    port map (
            in0 => \N__3416\,
            in1 => \N__3530\,
            in2 => \N__3556\,
            in3 => \N__3454\,
            lcout => pwm_cnte_0_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_togl_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__3443\,
            in1 => \N__3418\,
            in2 => \N__3535\,
            in3 => \N__3541\,
            lcout => \pwm_toglZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4391\,
            ce => 'H',
            sr => \N__4305\
        );

    \pwm_loc_RNO_1_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000100"
        )
    port map (
            in0 => \N__3397\,
            in1 => \N__3529\,
            in2 => \N__3448\,
            in3 => \N__3505\,
            lcout => OPEN,
            ltout => \pwm_loc_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pwm_loc_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110001010100"
        )
    port map (
            in0 => \N__3499\,
            in1 => \N__3480\,
            in2 => \N__3493\,
            in3 => \N__3417\,
            lcout => \pwm_locZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4391\,
            ce => 'H',
            sr => \N__4305\
        );

    \proc_pwm_fsm_pwm_loc20_0_I_33_c_RNIKR9E_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3440\,
            in2 => \_gnd_net_\,
            in3 => \N__3468\,
            lcout => \N_87\,
            ltout => \N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIVGJ71_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__3442\,
            in1 => \N__3415\,
            in2 => \N__3400\,
            in3 => \N__3396\,
            lcout => \N_78_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_RNO_0_0_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3321\,
            in2 => \_gnd_net_\,
            in3 => \N__3304\,
            lcout => prescale_cnt_s_0,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => prescale_cnt_cry_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3738\,
            in1 => \N__3657\,
            in2 => \_gnd_net_\,
            in3 => \N__3646\,
            lcout => \prescale_cntZ0Z_1\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_0,
            carryout => prescale_cnt_cry_1,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_2_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3731\,
            in1 => \N__4125\,
            in2 => \_gnd_net_\,
            in3 => \N__3643\,
            lcout => \prescale_cntZ0Z_2\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_1,
            carryout => prescale_cnt_cry_2,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_3_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3739\,
            in1 => \N__4149\,
            in2 => \_gnd_net_\,
            in3 => \N__3640\,
            lcout => \prescale_cntZ0Z_3\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_2,
            carryout => prescale_cnt_cry_3,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_4_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3732\,
            in1 => \N__4716\,
            in2 => \_gnd_net_\,
            in3 => \N__3637\,
            lcout => \prescale_cntZ0Z_4\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_3,
            carryout => prescale_cnt_cry_4,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_5_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3740\,
            in1 => \N__3864\,
            in2 => \_gnd_net_\,
            in3 => \N__3634\,
            lcout => \prescale_cntZ0Z_5\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_4,
            carryout => prescale_cnt_cry_5,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_6_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3733\,
            in1 => \N__3627\,
            in2 => \_gnd_net_\,
            in3 => \N__3616\,
            lcout => \prescale_cntZ0Z_6\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_5,
            carryout => prescale_cnt_cry_6,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_7_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3741\,
            in1 => \N__3609\,
            in2 => \_gnd_net_\,
            in3 => \N__3598\,
            lcout => \prescale_cntZ0Z_7\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_6,
            carryout => prescale_cnt_cry_7,
            clk => \N__4398\,
            ce => 'H',
            sr => \N__4311\
        );

    \prescale_cnt_8_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3730\,
            in1 => \N__3978\,
            in2 => \_gnd_net_\,
            in3 => \N__3595\,
            lcout => \prescale_cntZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => prescale_cnt_cry_8,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_9_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3737\,
            in1 => \N__3954\,
            in2 => \_gnd_net_\,
            in3 => \N__3793\,
            lcout => \prescale_cntZ0Z_9\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_8,
            carryout => prescale_cnt_cry_9,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_10_LC_3_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3727\,
            in1 => \N__3786\,
            in2 => \_gnd_net_\,
            in3 => \N__3775\,
            lcout => \prescale_cntZ0Z_10\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_9,
            carryout => prescale_cnt_cry_10,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_11_LC_3_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3734\,
            in1 => \N__3768\,
            in2 => \_gnd_net_\,
            in3 => \N__3757\,
            lcout => \prescale_cntZ0Z_11\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_10,
            carryout => prescale_cnt_cry_11,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_12_LC_3_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3728\,
            in1 => \N__4203\,
            in2 => \_gnd_net_\,
            in3 => \N__3754\,
            lcout => \prescale_cntZ0Z_12\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_11,
            carryout => prescale_cnt_cry_12,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_13_LC_3_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3735\,
            in1 => \N__4101\,
            in2 => \_gnd_net_\,
            in3 => \N__3751\,
            lcout => \prescale_cntZ0Z_13\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_12,
            carryout => prescale_cnt_cry_13,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_14_LC_3_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3729\,
            in1 => \N__3837\,
            in2 => \_gnd_net_\,
            in3 => \N__3748\,
            lcout => \prescale_cntZ0Z_14\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_13,
            carryout => prescale_cnt_cry_14,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_15_LC_3_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3736\,
            in1 => \N__3810\,
            in2 => \_gnd_net_\,
            in3 => \N__3745\,
            lcout => \prescale_cntZ0Z_15\,
            ltout => OPEN,
            carryin => prescale_cnt_cry_14,
            carryout => prescale_cnt_cry_15,
            clk => \N__4399\,
            ce => 'H',
            sr => \N__4315\
        );

    \prescale_cnt_16_LC_3_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__3742\,
            in1 => \N__4188\,
            in2 => \_gnd_net_\,
            in3 => \N__3679\,
            lcout => \prescale_cntZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4403\,
            ce => 'H',
            sr => \N__4320\
        );

    \prescale_stop_p1_0_LC_3_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4678\,
            in1 => \N__4597\,
            in2 => \_gnd_net_\,
            in3 => \N__4461\,
            lcout => \prescale_stop_p1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4403\,
            ce => 'H',
            sr => \N__4320\
        );

    \prescale_stop_p1_1_LC_3_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__4462\,
            in1 => \N__4598\,
            in2 => \_gnd_net_\,
            in3 => \N__4679\,
            lcout => \prescale_stop_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4403\,
            ce => 'H',
            sr => \N__4320\
        );

    \pwm_lout_p1_4_LC_3_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3898\,
            lcout => \pwm_lout_p1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4408\,
            ce => 'H',
            sr => \N__4327\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_15_c_RNO_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__4227\,
            in1 => \N__3799\,
            in2 => \N__3853\,
            in3 => \N__3826\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_p1_5_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3871\,
            lcout => \prescale_cnt_p1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4400\,
            ce => 'H',
            sr => \N__4324\
        );

    \prescale_stop_p1_14_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4687\,
            in1 => \N__4573\,
            in2 => \_gnd_net_\,
            in3 => \N__4489\,
            lcout => \prescale_stop_p1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4400\,
            ce => 'H',
            sr => \N__4324\
        );

    \prescale_stop_p1_15_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4162\,
            lcout => \prescale_stop_p1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4400\,
            ce => 'H',
            sr => \N__4324\
        );

    \prescale_cnt_p1_14_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3844\,
            lcout => \prescale_cnt_p1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4400\,
            ce => 'H',
            sr => \N__4324\
        );

    \prescale_cnt_p1_15_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3820\,
            lcout => \prescale_cnt_p1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4400\,
            ce => 'H',
            sr => \N__4324\
        );

    \prescale_stop_p1_8_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4688\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \prescale_stop_p1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4392\,
            ce => 'H',
            sr => \N__4321\
        );

    \prescale_stop_p1_2_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4689\,
            lcout => \prescale_stop_p1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4392\,
            ce => 'H',
            sr => \N__4321\
        );

    \pwm_prescale_p1_1_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \pwm_prescale_p1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4392\,
            ce => 'H',
            sr => \N__4321\
        );

    \pwm_lout_p1_5_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4021\,
            lcout => \pwm_lout_p1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4392\,
            ce => 'H',
            sr => \N__4321\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_33_c_RNO_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3943\,
            in1 => \N__3967\,
            in2 => \N__3994\,
            in3 => \N__3937\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_p1_8_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3985\,
            lcout => \prescale_cnt_p1Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4401\,
            ce => 'H',
            sr => \N__4312\
        );

    \prescale_cnt_p1_9_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3961\,
            lcout => \prescale_cnt_p1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4401\,
            ce => 'H',
            sr => \N__4312\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_51_c_RNO_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__3936\,
            in1 => \N__4138\,
            in2 => \N__3928\,
            in3 => \N__4114\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_stop_p1_3_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4698\,
            in1 => \N__4575\,
            in2 => \_gnd_net_\,
            in3 => \N__4478\,
            lcout => \prescale_stop_p1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4401\,
            ce => 'H',
            sr => \N__4312\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_1_c_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3919\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_0,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_51_c_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4090\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_0,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_45_c_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4237\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_1,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_39_c_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4084\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_2,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_33_c_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4072\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_3,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_27_c_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4066\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_4,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_21_c_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4504\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_5,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_15_c_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4054\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => proc_pwm_cnt_prescale_cnt10_0_data_tmp_6,
            carryout => proc_pwm_cnt_prescale_cnt10_0_data_tmp_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_9_c_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4216\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => proc_pwm_cnt_prescale_cnt10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_THRU_LUT4_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4045\,
            lcout => \proc_pwm_cnt_prescale_cnt10_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_45_c_RNO_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__4728\,
            in1 => \N__4705\,
            in2 => \N__4171\,
            in3 => \N__4246\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNO_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__4177\,
            in1 => \N__4729\,
            in2 => \_gnd_net_\,
            in3 => \N__4231\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_p1_12_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4210\,
            lcout => \prescale_cnt_p1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => 'H',
            sr => \N__4325\
        );

    \prescale_cnt_p1_16_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4192\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \prescale_cnt_p1Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => 'H',
            sr => \N__4325\
        );

    \prescale_stop_p1_5_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000100010"
        )
    port map (
            in0 => \N__4699\,
            in1 => \N__4595\,
            in2 => \_gnd_net_\,
            in3 => \N__4479\,
            lcout => \prescale_stop_p1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4406\,
            ce => 'H',
            sr => \N__4325\
        );

    \prescale_stop_1_8_3__m8_0_a3_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4680\,
            in2 => \_gnd_net_\,
            in3 => \N__4488\,
            lcout => prescale_stop_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_cnt_p1_3_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4156\,
            lcout => \prescale_cnt_p1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4402\,
            ce => 'H',
            sr => \N__4316\
        );

    \prescale_cnt_p1_2_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4132\,
            lcout => \prescale_cnt_p1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4402\,
            ce => 'H',
            sr => \N__4316\
        );

    \prescale_cnt_p1_13_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4108\,
            lcout => \prescale_cnt_p1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4402\,
            ce => 'H',
            sr => \N__4316\
        );

    \prescale_stop_p1_4_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4594\,
            in2 => \_gnd_net_\,
            in3 => \N__4697\,
            lcout => \prescale_stop_p1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4404\,
            ce => 'H',
            sr => \N__4322\
        );

    \prescale_cnt_p1_4_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4720\,
            lcout => \prescale_cnt_p1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4404\,
            ce => 'H',
            sr => \N__4322\
        );

    \prescale_stop_1_8_3__m4_0_a3_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4696\,
            in2 => \_gnd_net_\,
            in3 => \N__4593\,
            lcout => prescale_stop_1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \proc_pwm_cnt_prescale_cnt10_0_I_21_c_RNO_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__4414\,
            in1 => \N__4519\,
            in2 => \_gnd_net_\,
            in3 => \N__4510\,
            lcout => \proc_pwm_cnt_prescale_cnt10_0_N_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \prescale_stop_p1_13_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4498\,
            in2 => \_gnd_net_\,
            in3 => \N__4480\,
            lcout => \prescale_stop_p1Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4407\,
            ce => 'H',
            sr => \N__4326\
        );
end \INTERFACE\;
