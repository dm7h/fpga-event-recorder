// ******************************************************************************

// iCEcube Netlister

// Version:            2015.04.27409

// Build Date:         May 27 2015 16:13:33

// File Generated:     Feb 6 2017 16:52:10

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "gpio_pwm" view "INTERFACE"

module gpio_pwm (
    pwm_prescale,
    pwm_ctrl,
    pwm_hout,
    pwm_lout,
    clk,
    pwm_pin,
    reset);

    input [2:0] pwm_prescale;
    input [1:0] pwm_ctrl;
    input [11:0] pwm_hout;
    input [11:0] pwm_lout;
    input clk;
    output pwm_pin;
    input reset;

    wire N__5030;
    wire N__5029;
    wire N__5028;
    wire N__5020;
    wire N__5019;
    wire N__5018;
    wire N__5009;
    wire N__5008;
    wire N__5007;
    wire N__5000;
    wire N__4999;
    wire N__4998;
    wire N__4991;
    wire N__4990;
    wire N__4989;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4973;
    wire N__4972;
    wire N__4971;
    wire N__4964;
    wire N__4963;
    wire N__4962;
    wire N__4955;
    wire N__4954;
    wire N__4953;
    wire N__4946;
    wire N__4945;
    wire N__4944;
    wire N__4937;
    wire N__4936;
    wire N__4935;
    wire N__4928;
    wire N__4927;
    wire N__4926;
    wire N__4919;
    wire N__4918;
    wire N__4917;
    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4901;
    wire N__4900;
    wire N__4899;
    wire N__4892;
    wire N__4891;
    wire N__4890;
    wire N__4883;
    wire N__4882;
    wire N__4881;
    wire N__4874;
    wire N__4873;
    wire N__4872;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4856;
    wire N__4855;
    wire N__4854;
    wire N__4847;
    wire N__4846;
    wire N__4845;
    wire N__4838;
    wire N__4837;
    wire N__4836;
    wire N__4829;
    wire N__4828;
    wire N__4827;
    wire N__4820;
    wire N__4819;
    wire N__4818;
    wire N__4811;
    wire N__4810;
    wire N__4809;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4793;
    wire N__4792;
    wire N__4791;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4766;
    wire N__4765;
    wire N__4764;
    wire N__4757;
    wire N__4756;
    wire N__4755;
    wire N__4748;
    wire N__4747;
    wire N__4746;
    wire N__4729;
    wire N__4728;
    wire N__4723;
    wire N__4720;
    wire N__4717;
    wire N__4716;
    wire N__4713;
    wire N__4710;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4698;
    wire N__4697;
    wire N__4696;
    wire N__4693;
    wire N__4690;
    wire N__4689;
    wire N__4688;
    wire N__4687;
    wire N__4684;
    wire N__4681;
    wire N__4680;
    wire N__4679;
    wire N__4678;
    wire N__4673;
    wire N__4668;
    wire N__4667;
    wire N__4666;
    wire N__4665;
    wire N__4662;
    wire N__4657;
    wire N__4654;
    wire N__4649;
    wire N__4648;
    wire N__4643;
    wire N__4636;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4615;
    wire N__4610;
    wire N__4603;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4597;
    wire N__4596;
    wire N__4595;
    wire N__4594;
    wire N__4593;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4579;
    wire N__4576;
    wire N__4575;
    wire N__4574;
    wire N__4573;
    wire N__4572;
    wire N__4569;
    wire N__4566;
    wire N__4563;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4545;
    wire N__4542;
    wire N__4537;
    wire N__4532;
    wire N__4519;
    wire N__4516;
    wire N__4513;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4498;
    wire N__4495;
    wire N__4492;
    wire N__4491;
    wire N__4490;
    wire N__4489;
    wire N__4488;
    wire N__4481;
    wire N__4480;
    wire N__4479;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4453;
    wire N__4450;
    wire N__4445;
    wire N__4440;
    wire N__4435;
    wire N__4434;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4414;
    wire N__4411;
    wire N__4408;
    wire N__4407;
    wire N__4406;
    wire N__4405;
    wire N__4404;
    wire N__4403;
    wire N__4402;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4397;
    wire N__4396;
    wire N__4395;
    wire N__4394;
    wire N__4393;
    wire N__4392;
    wire N__4391;
    wire N__4390;
    wire N__4389;
    wire N__4388;
    wire N__4387;
    wire N__4386;
    wire N__4385;
    wire N__4384;
    wire N__4333;
    wire N__4330;
    wire N__4327;
    wire N__4326;
    wire N__4325;
    wire N__4324;
    wire N__4323;
    wire N__4322;
    wire N__4321;
    wire N__4320;
    wire N__4319;
    wire N__4318;
    wire N__4317;
    wire N__4316;
    wire N__4315;
    wire N__4314;
    wire N__4313;
    wire N__4312;
    wire N__4311;
    wire N__4310;
    wire N__4309;
    wire N__4308;
    wire N__4307;
    wire N__4306;
    wire N__4305;
    wire N__4304;
    wire N__4303;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4237;
    wire N__4234;
    wire N__4231;
    wire N__4228;
    wire N__4227;
    wire N__4224;
    wire N__4221;
    wire N__4216;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4203;
    wire N__4200;
    wire N__4197;
    wire N__4192;
    wire N__4189;
    wire N__4188;
    wire N__4185;
    wire N__4182;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4149;
    wire N__4146;
    wire N__4143;
    wire N__4138;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4125;
    wire N__4122;
    wire N__4119;
    wire N__4114;
    wire N__4111;
    wire N__4108;
    wire N__4105;
    wire N__4102;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4090;
    wire N__4087;
    wire N__4084;
    wire N__4081;
    wire N__4078;
    wire N__4075;
    wire N__4072;
    wire N__4069;
    wire N__4066;
    wire N__4063;
    wire N__4060;
    wire N__4057;
    wire N__4054;
    wire N__4051;
    wire N__4048;
    wire N__4045;
    wire N__4042;
    wire N__4041;
    wire N__4036;
    wire N__4033;
    wire N__4030;
    wire N__4027;
    wire N__4024;
    wire N__4021;
    wire N__4018;
    wire N__4015;
    wire N__4012;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3997;
    wire N__3994;
    wire N__3991;
    wire N__3988;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3967;
    wire N__3964;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3954;
    wire N__3951;
    wire N__3948;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3936;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3889;
    wire N__3886;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3865;
    wire N__3864;
    wire N__3861;
    wire N__3858;
    wire N__3853;
    wire N__3850;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3837;
    wire N__3834;
    wire N__3831;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3799;
    wire N__3796;
    wire N__3793;
    wire N__3790;
    wire N__3787;
    wire N__3786;
    wire N__3783;
    wire N__3780;
    wire N__3775;
    wire N__3772;
    wire N__3769;
    wire N__3768;
    wire N__3765;
    wire N__3762;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3741;
    wire N__3740;
    wire N__3739;
    wire N__3738;
    wire N__3737;
    wire N__3736;
    wire N__3735;
    wire N__3734;
    wire N__3733;
    wire N__3732;
    wire N__3731;
    wire N__3730;
    wire N__3729;
    wire N__3728;
    wire N__3727;
    wire N__3724;
    wire N__3715;
    wire N__3706;
    wire N__3699;
    wire N__3690;
    wire N__3679;
    wire N__3676;
    wire N__3675;
    wire N__3674;
    wire N__3673;
    wire N__3668;
    wire N__3663;
    wire N__3658;
    wire N__3657;
    wire N__3654;
    wire N__3651;
    wire N__3646;
    wire N__3643;
    wire N__3640;
    wire N__3637;
    wire N__3634;
    wire N__3631;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3609;
    wire N__3606;
    wire N__3603;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3591;
    wire N__3588;
    wire N__3585;
    wire N__3580;
    wire N__3577;
    wire N__3576;
    wire N__3573;
    wire N__3570;
    wire N__3567;
    wire N__3564;
    wire N__3559;
    wire N__3556;
    wire N__3553;
    wire N__3552;
    wire N__3549;
    wire N__3546;
    wire N__3541;
    wire N__3538;
    wire N__3535;
    wire N__3534;
    wire N__3531;
    wire N__3530;
    wire N__3529;
    wire N__3526;
    wire N__3519;
    wire N__3516;
    wire N__3513;
    wire N__3510;
    wire N__3505;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3480;
    wire N__3477;
    wire N__3474;
    wire N__3469;
    wire N__3468;
    wire N__3467;
    wire N__3464;
    wire N__3459;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3444;
    wire N__3443;
    wire N__3442;
    wire N__3441;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3425;
    wire N__3418;
    wire N__3417;
    wire N__3416;
    wire N__3415;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3396;
    wire N__3395;
    wire N__3388;
    wire N__3387;
    wire N__3384;
    wire N__3381;
    wire N__3378;
    wire N__3373;
    wire N__3372;
    wire N__3371;
    wire N__3370;
    wire N__3369;
    wire N__3368;
    wire N__3359;
    wire N__3358;
    wire N__3357;
    wire N__3356;
    wire N__3355;
    wire N__3354;
    wire N__3353;
    wire N__3348;
    wire N__3345;
    wire N__3340;
    wire N__3331;
    wire N__3322;
    wire N__3321;
    wire N__3318;
    wire N__3315;
    wire N__3310;
    wire N__3307;
    wire N__3304;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3283;
    wire N__3280;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3255;
    wire N__3254;
    wire N__3251;
    wire N__3248;
    wire N__3245;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3228;
    wire N__3225;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3208;
    wire N__3205;
    wire N__3202;
    wire N__3199;
    wire N__3196;
    wire N__3193;
    wire N__3192;
    wire N__3189;
    wire N__3188;
    wire N__3185;
    wire N__3182;
    wire N__3179;
    wire N__3172;
    wire N__3171;
    wire N__3170;
    wire N__3167;
    wire N__3164;
    wire N__3161;
    wire N__3154;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3142;
    wire N__3139;
    wire N__3136;
    wire N__3133;
    wire N__3130;
    wire N__3127;
    wire N__3124;
    wire N__3121;
    wire N__3118;
    wire N__3115;
    wire N__3112;
    wire N__3109;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3094;
    wire N__3091;
    wire N__3088;
    wire N__3085;
    wire N__3082;
    wire N__3079;
    wire N__3076;
    wire N__3073;
    wire N__3070;
    wire N__3067;
    wire N__3064;
    wire N__3061;
    wire N__3058;
    wire N__3055;
    wire N__3052;
    wire N__3049;
    wire N__3046;
    wire N__3043;
    wire N__3040;
    wire N__3037;
    wire N__3034;
    wire N__3033;
    wire N__3032;
    wire N__3025;
    wire N__3022;
    wire N__3021;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3001;
    wire N__3000;
    wire N__2999;
    wire N__2996;
    wire N__2993;
    wire N__2990;
    wire N__2987;
    wire N__2980;
    wire N__2977;
    wire N__2974;
    wire N__2971;
    wire N__2968;
    wire N__2967;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2950;
    wire N__2947;
    wire N__2946;
    wire N__2945;
    wire N__2942;
    wire N__2937;
    wire N__2932;
    wire N__2929;
    wire N__2926;
    wire N__2923;
    wire N__2922;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2905;
    wire N__2902;
    wire N__2901;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2884;
    wire N__2881;
    wire N__2880;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2860;
    wire N__2857;
    wire N__2856;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire N__2846;
    wire N__2843;
    wire N__2836;
    wire N__2833;
    wire N__2830;
    wire N__2827;
    wire N__2824;
    wire N__2821;
    wire N__2818;
    wire N__2815;
    wire N__2812;
    wire N__2809;
    wire N__2806;
    wire N__2803;
    wire N__2800;
    wire N__2797;
    wire N__2794;
    wire N__2791;
    wire N__2788;
    wire N__2785;
    wire N__2782;
    wire N__2779;
    wire N__2776;
    wire N__2773;
    wire N__2770;
    wire N__2767;
    wire N__2764;
    wire N__2761;
    wire N__2758;
    wire N__2755;
    wire N__2752;
    wire N__2749;
    wire N__2746;
    wire N__2743;
    wire N__2740;
    wire N__2737;
    wire N__2734;
    wire N__2731;
    wire N__2728;
    wire N__2725;
    wire N__2722;
    wire N__2719;
    wire N__2716;
    wire N__2713;
    wire N__2710;
    wire N__2707;
    wire N__2704;
    wire N__2701;
    wire N__2698;
    wire N__2695;
    wire N__2692;
    wire N__2689;
    wire N__2686;
    wire N__2683;
    wire N__2680;
    wire N__2677;
    wire N__2674;
    wire N__2671;
    wire N__2668;
    wire N__2665;
    wire N__2662;
    wire N__2659;
    wire N__2656;
    wire N__2653;
    wire N__2650;
    wire N__2647;
    wire N__2644;
    wire N__2641;
    wire N__2638;
    wire N__2635;
    wire N__2632;
    wire N__2629;
    wire N__2626;
    wire N__2623;
    wire N__2620;
    wire N__2617;
    wire N__2614;
    wire N__2611;
    wire N__2608;
    wire N__2605;
    wire N__2602;
    wire N__2599;
    wire N__2596;
    wire N__2593;
    wire N__2590;
    wire N__2587;
    wire N__2584;
    wire N__2581;
    wire N__2578;
    wire N__2575;
    wire N__2572;
    wire N__2569;
    wire N__2566;
    wire N__2563;
    wire N__2560;
    wire N__2557;
    wire N__2554;
    wire N__2551;
    wire N__2548;
    wire N__2545;
    wire N__2542;
    wire N__2539;
    wire N__2536;
    wire N__2533;
    wire N__2530;
    wire N__2527;
    wire N__2524;
    wire N__2521;
    wire N__2518;
    wire N__2515;
    wire N__2512;
    wire N__2509;
    wire N__2506;
    wire N__2503;
    wire N__2500;
    wire N__2497;
    wire N__2494;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2482;
    wire N__2479;
    wire N__2476;
    wire N__2473;
    wire N__2470;
    wire N__2467;
    wire N__2464;
    wire N__2461;
    wire N__2458;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2437;
    wire N__2434;
    wire N__2431;
    wire N__2428;
    wire N__2425;
    wire N__2422;
    wire N__2419;
    wire N__2416;
    wire N__2413;
    wire N__2410;
    wire N__2407;
    wire N__2404;
    wire N__2401;
    wire N__2398;
    wire N__2395;
    wire N__2392;
    wire N__2389;
    wire N__2386;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2374;
    wire N__2371;
    wire N__2368;
    wire N__2365;
    wire N__2362;
    wire N__2359;
    wire N__2356;
    wire N__2353;
    wire N__2350;
    wire N__2347;
    wire N__2344;
    wire N__2341;
    wire N__2338;
    wire N__2335;
    wire N__2332;
    wire N__2329;
    wire N__2326;
    wire N__2323;
    wire N__2320;
    wire N__2317;
    wire N__2314;
    wire N__2311;
    wire N__2308;
    wire N__2305;
    wire N__2302;
    wire N__2299;
    wire N__2296;
    wire N__2293;
    wire N__2290;
    wire N__2287;
    wire N__2284;
    wire N__2281;
    wire N__2278;
    wire N__2275;
    wire N__2272;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire VCCG0;
    wire GNDG0;
    wire pwm_pin_c;
    wire pwm_lout_c_9;
    wire pwm_lout_c_6;
    wire pwm_hout_c_9;
    wire pwm_hout_c_8;
    wire bfn_1_10_0_;
    wire proc_pwm_fsm_pwm_loc8_0_data_tmp_0;
    wire proc_pwm_fsm_pwm_loc8_0_data_tmp_1;
    wire proc_pwm_fsm_pwm_loc8_0_data_tmp_2;
    wire proc_pwm_fsm_pwm_loc8_0_data_tmp_3;
    wire proc_pwm_fsm_pwm_loc8_0_data_tmp_4;
    wire proc_pwm_fsm_pwm_loc8;
    wire pwm_lout_p1Z0Z_6;
    wire proc_pwm_fsm_pwm_loc8_0_N_26;
    wire proc_pwm_fsm_pwm_loc8_0_N_6;
    wire proc_pwm_fsm_pwm_loc8_0_N_16;
    wire proc_pwm_fsm_pwm_loc8_0_N_21;
    wire pwm_hout_p1Z0Z_8;
    wire pwm_hout_p1Z0Z_9;
    wire proc_pwm_fsm_pwm_loc8_0_N_11;
    wire pwm_hout_c_5;
    wire pwm_hout_p1Z0Z_5;
    wire pwm_hout_c_4;
    wire pwm_hout_p1Z0Z_4;
    wire pwm_hout_c_0;
    wire pwm_hout_p1Z0Z_0;
    wire pwm_hout_c_3;
    wire pwm_hout_p1Z0Z_3;
    wire pwm_lout_c_2;
    wire pwm_lout_p1Z0Z_2;
    wire pwm_hout_c_1;
    wire pwm_hout_p1Z0Z_1;
    wire pwm_hout_c_2;
    wire pwm_hout_p1Z0Z_2;
    wire pwm_lout_c_3;
    wire pwm_lout_p1Z0Z_3;
    wire proc_pwm_fsm_pwm_loc8_0_N_1;
    wire pwm_hout_c_6;
    wire pwm_hout_p1Z0Z_6;
    wire pwm_hout_c_10;
    wire pwm_hout_p1Z0Z_10;
    wire pwm_hout_c_7;
    wire pwm_hout_p1Z0Z_7;
    wire pwm_hout_c_11;
    wire pwm_hout_p1Z0Z_11;
    wire pwm_prescale_c_0;
    wire pwm_lout_c_7;
    wire pwm_lout_p1Z0Z_7;
    wire pwm_prescale_c_2;
    wire pwm_lout_c_8;
    wire pwm_ctrl_c_0;
    wire pwm_lout_p1Z0Z_8;
    wire pwm_lout_p1Z0Z_9;
    wire bfn_2_10_0_;
    wire proc_pwm_fsm_pwm_loc20_0_N_21;
    wire proc_pwm_fsm_pwm_loc20_0_data_tmp_0;
    wire proc_pwm_fsm_pwm_loc20_0_data_tmp_1;
    wire proc_pwm_fsm_pwm_loc20_0_N_6;
    wire proc_pwm_fsm_pwm_loc20_0_data_tmp_2;
    wire proc_pwm_fsm_pwm_loc20_0_N_11;
    wire proc_pwm_fsm_pwm_loc20_0_data_tmp_3;
    wire proc_pwm_fsm_pwm_loc20_0_data_tmp_4;
    wire proc_pwm_fsm_pwm_loc20;
    wire bfn_2_11_0_;
    wire pwm_cnt_cry_0;
    wire pwm_cntZ0Z_2;
    wire pwm_cnt_cry_1;
    wire pwm_cntZ0Z_3;
    wire pwm_cnt_cry_2;
    wire pwm_cnt_cry_3;
    wire pwm_cnt_cry_4;
    wire pwm_cntZ0Z_6;
    wire pwm_cnt_cry_5;
    wire pwm_cntZ0Z_7;
    wire pwm_cnt_cry_6;
    wire pwm_cnt_cry_7;
    wire pwm_cntZ0Z_8;
    wire bfn_2_12_0_;
    wire pwm_cntZ0Z_9;
    wire pwm_cnt_cry_8;
    wire pwm_cnt_cry_9;
    wire pwm_cnt_cry_10;
    wire N_8_cascade_;
    wire prescale_cnt_p1Z0Z_0;
    wire prescale_cnt_p1Z0Z_1;
    wire N_38;
    wire pwm_cntZ0Z_11;
    wire pwm_cntZ0Z_10;
    wire proc_pwm_fsm_pwm_loc20_0_N_1;
    wire pwm_lout_c_11;
    wire pwm_lout_p1Z0Z_11;
    wire pwm_lout_c_10;
    wire pwm_lout_p1Z0Z_10;
    wire pwm_lout_c_1;
    wire pwm_ctrl_c_1;
    wire pwm_lout_c_0;
    wire prescale_stop_p1Z0Z_6;
    wire prescale_cnt_p1Z0Z_7;
    wire prescale_stop_p1Z0Z_7;
    wire prescale_cnt_p1Z0Z_6;
    wire prescale_stop_p1Z0Z_10;
    wire prescale_cnt_p1Z0Z_11;
    wire prescale_cnt_p1Z0Z_10;
    wire pwm_cntZ0Z_1;
    wire pwm_lout_p1Z0Z_1;
    wire pwm_cntZ0Z_0;
    wire pwm_lout_p1Z0Z_0;
    wire proc_pwm_fsm_pwm_loc20_0_N_26;
    wire pwm_cntZ0Z_5;
    wire pwm_cntZ0Z_4;
    wire proc_pwm_fsm_pwm_loc20_0_N_16;
    wire pwm_ctrl_p1Z0Z_0;
    wire pwm_ctrl_p1Z0Z_1;
    wire pwm_loc_1_sqmuxa_cascade_;
    wire un1_pwm_loc8_1_0_cascade_;
    wire pwm_cnte_0_i;
    wire un1_pwm_loc8_1_0;
    wire prescale_tickZ0;
    wire pwm_loc_1_sqmuxa;
    wire pwm_loc_0_sqmuxa_1;
    wire pwm_loc_1_sqmuxa_1_cascade_;
    wire pwm_locZ0;
    wire proc_pwm_fsm_pwm_loc20_THRU_CO;
    wire N_87;
    wire pwm_toglZ0;
    wire N_86;
    wire N_87_cascade_;
    wire proc_pwm_fsm_pwm_loc8_THRU_CO;
    wire N_78_0_i;
    wire prescale_cntZ0Z_0;
    wire prescale_cnt_s_0;
    wire bfn_3_12_0_;
    wire prescale_cntZ0Z_1;
    wire prescale_cnt_cry_0;
    wire prescale_cnt_cry_1;
    wire prescale_cnt_cry_2;
    wire prescale_cnt_cry_3;
    wire prescale_cnt_cry_4;
    wire prescale_cntZ0Z_6;
    wire prescale_cnt_cry_5;
    wire prescale_cntZ0Z_7;
    wire prescale_cnt_cry_6;
    wire prescale_cnt_cry_7;
    wire bfn_3_13_0_;
    wire prescale_cnt_cry_8;
    wire prescale_cntZ0Z_10;
    wire prescale_cnt_cry_9;
    wire prescale_cntZ0Z_11;
    wire prescale_cnt_cry_10;
    wire prescale_cnt_cry_11;
    wire prescale_cnt_cry_12;
    wire prescale_cnt_cry_13;
    wire prescale_cnt_cry_14;
    wire prescale_cnt_cry_15;
    wire N_8;
    wire bfn_3_14_0_;
    wire prescale_stop_p1Z0Z_0;
    wire prescale_stop_p1Z0Z_1;
    wire pwm_lout_c_4;
    wire pwm_lout_p1Z0Z_4;
    wire prescale_cntZ0Z_5;
    wire prescale_stop_p1Z0Z_15;
    wire prescale_cntZ0Z_14;
    wire prescale_cnt_p1Z0Z_14;
    wire prescale_cntZ0Z_15;
    wire prescale_cnt_p1Z0Z_15;
    wire pwm_prescale_c_1;
    wire pwm_lout_c_5;
    wire pwm_lout_p1Z0Z_5;
    wire prescale_stop_p1Z0Z_8;
    wire prescale_cntZ0Z_8;
    wire prescale_cnt_p1Z0Z_8;
    wire prescale_cntZ0Z_9;
    wire prescale_cnt_p1Z0Z_9;
    wire prescale_stop_p1Z0Z_2;
    wire prescale_stop_p1Z0Z_3;
    wire proc_pwm_cnt_prescale_cnt10_0_N_41;
    wire bfn_5_12_0_;
    wire proc_pwm_cnt_prescale_cnt10_0_N_1;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_0;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_1;
    wire proc_pwm_cnt_prescale_cnt10_0_N_11;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_2;
    wire proc_pwm_cnt_prescale_cnt10_0_N_16;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_3;
    wire proc_pwm_cnt_prescale_cnt10_0_N_21;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_4;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_5;
    wire proc_pwm_cnt_prescale_cnt10_0_N_31;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_6;
    wire proc_pwm_cnt_prescale_cnt10_0_data_tmp_7;
    wire bfn_5_13_0_;
    wire proc_pwm_cnt_prescale_cnt10;
    wire proc_pwm_cnt_prescale_cnt10_THRU_CO;
    wire prescale_cnt_p1Z0Z_5;
    wire proc_pwm_cnt_prescale_cnt10_0_N_6;
    wire prescale_stop_p1Z0Z_14;
    wire proc_pwm_cnt_prescale_cnt10_0_N_36;
    wire prescale_cntZ0Z_12;
    wire prescale_cntZ0Z_16;
    wire prescale_cnt_p1Z0Z_16;
    wire prescale_stop_p1Z0Z_5;
    wire prescale_stop_1_7;
    wire prescale_cntZ0Z_3;
    wire prescale_cnt_p1Z0Z_3;
    wire prescale_cntZ0Z_2;
    wire prescale_cnt_p1Z0Z_2;
    wire prescale_cntZ0Z_13;
    wire prescale_stop_p1Z0Z_4;
    wire prescale_cntZ0Z_4;
    wire prescale_cnt_p1Z0Z_4;
    wire pwm_prescale_p1Z0Z_2;
    wire pwm_prescale_p1Z0Z_1;
    wire prescale_cnt_p1Z0Z_13;
    wire prescale_cnt_p1Z0Z_12;
    wire proc_pwm_cnt_prescale_cnt10_0_N_26;
    wire prescale_stop_1_8;
    wire pwm_prescale_p1Z0Z_0;
    wire prescale_stop_p1Z0Z_13;
    wire _gnd_net_;
    wire clk_c_g;
    wire reset_c_g;

    PRE_IO_GBUF reset_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5028),
            .GLOBALBUFFEROUTPUT(reset_c_g));
    IO_PAD reset_ibuf_gb_io_iopad (
            .OE(N__5030),
            .DIN(N__5029),
            .DOUT(N__5028),
            .PACKAGEPIN(reset));
    defparam reset_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam reset_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO reset_ibuf_gb_io_preio (
            .PADOEN(N__5030),
            .PADOUT(N__5029),
            .PADIN(N__5028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    PRE_IO_GBUF clk_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__5018),
            .GLOBALBUFFEROUTPUT(clk_c_g));
    IO_PAD clk_ibuf_gb_io_iopad (
            .OE(N__5020),
            .DIN(N__5019),
            .DOUT(N__5018),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_gb_io_preio (
            .PADOEN(N__5020),
            .PADOUT(N__5019),
            .PADIN(N__5018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_11_iopad (
            .OE(N__5009),
            .DIN(N__5008),
            .DOUT(N__5007),
            .PACKAGEPIN(pwm_hout[11]));
    defparam pwm_hout_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_11_preio (
            .PADOEN(N__5009),
            .PADOUT(N__5008),
            .PADIN(N__5007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_5_iopad (
            .OE(N__5000),
            .DIN(N__4999),
            .DOUT(N__4998),
            .PACKAGEPIN(pwm_hout[5]));
    defparam pwm_hout_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_5_preio (
            .PADOEN(N__5000),
            .PADOUT(N__4999),
            .PADIN(N__4998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_2_iopad (
            .OE(N__4991),
            .DIN(N__4990),
            .DOUT(N__4989),
            .PACKAGEPIN(pwm_hout[2]));
    defparam pwm_hout_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_2_preio (
            .PADOEN(N__4991),
            .PADOUT(N__4990),
            .PADIN(N__4989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_4_iopad (
            .OE(N__4982),
            .DIN(N__4981),
            .DOUT(N__4980),
            .PACKAGEPIN(pwm_lout[4]));
    defparam pwm_lout_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_4_preio (
            .PADOEN(N__4982),
            .PADOUT(N__4981),
            .PADIN(N__4980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_ctrl_ibuf_0_iopad (
            .OE(N__4973),
            .DIN(N__4972),
            .DOUT(N__4971),
            .PACKAGEPIN(pwm_ctrl[0]));
    defparam pwm_ctrl_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam pwm_ctrl_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_ctrl_ibuf_0_preio (
            .PADOEN(N__4973),
            .PADOUT(N__4972),
            .PADIN(N__4971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_ctrl_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_9_iopad (
            .OE(N__4964),
            .DIN(N__4963),
            .DOUT(N__4962),
            .PACKAGEPIN(pwm_lout[9]));
    defparam pwm_lout_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_9_preio (
            .PADOEN(N__4964),
            .PADOUT(N__4963),
            .PADIN(N__4962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_prescale_ibuf_1_iopad (
            .OE(N__4955),
            .DIN(N__4954),
            .DOUT(N__4953),
            .PACKAGEPIN(pwm_prescale[1]));
    defparam pwm_prescale_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam pwm_prescale_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_prescale_ibuf_1_preio (
            .PADOEN(N__4955),
            .PADOUT(N__4954),
            .PADIN(N__4953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_prescale_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_7_iopad (
            .OE(N__4946),
            .DIN(N__4945),
            .DOUT(N__4944),
            .PACKAGEPIN(pwm_hout[7]));
    defparam pwm_hout_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_7_preio (
            .PADOEN(N__4946),
            .PADOUT(N__4945),
            .PADIN(N__4944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_1_iopad (
            .OE(N__4937),
            .DIN(N__4936),
            .DOUT(N__4935),
            .PACKAGEPIN(pwm_lout[1]));
    defparam pwm_lout_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_1_preio (
            .PADOEN(N__4937),
            .PADOUT(N__4936),
            .PADIN(N__4935),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_pin_obuf_iopad (
            .OE(N__4928),
            .DIN(N__4927),
            .DOUT(N__4926),
            .PACKAGEPIN(pwm_pin));
    defparam pwm_pin_obuf_preio.NEG_TRIGGER=1'b0;
    defparam pwm_pin_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO pwm_pin_obuf_preio (
            .PADOEN(N__4928),
            .PADOUT(N__4927),
            .PADIN(N__4926),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__2299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_6_iopad (
            .OE(N__4919),
            .DIN(N__4918),
            .DOUT(N__4917),
            .PACKAGEPIN(pwm_lout[6]));
    defparam pwm_lout_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_6_preio (
            .PADOEN(N__4919),
            .PADOUT(N__4918),
            .PADIN(N__4917),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_9_iopad (
            .OE(N__4910),
            .DIN(N__4909),
            .DOUT(N__4908),
            .PACKAGEPIN(pwm_hout[9]));
    defparam pwm_hout_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_9_preio (
            .PADOEN(N__4910),
            .PADOUT(N__4909),
            .PADIN(N__4908),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_4_iopad (
            .OE(N__4901),
            .DIN(N__4900),
            .DOUT(N__4899),
            .PACKAGEPIN(pwm_hout[4]));
    defparam pwm_hout_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_4_preio (
            .PADOEN(N__4901),
            .PADOUT(N__4900),
            .PADIN(N__4899),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_1_iopad (
            .OE(N__4892),
            .DIN(N__4891),
            .DOUT(N__4890),
            .PACKAGEPIN(pwm_hout[1]));
    defparam pwm_hout_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_1_preio (
            .PADOEN(N__4892),
            .PADOUT(N__4891),
            .PADIN(N__4890),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_3_iopad (
            .OE(N__4883),
            .DIN(N__4882),
            .DOUT(N__4881),
            .PACKAGEPIN(pwm_lout[3]));
    defparam pwm_lout_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_3_preio (
            .PADOEN(N__4883),
            .PADOUT(N__4882),
            .PADIN(N__4881),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_ctrl_ibuf_1_iopad (
            .OE(N__4874),
            .DIN(N__4873),
            .DOUT(N__4872),
            .PACKAGEPIN(pwm_ctrl[1]));
    defparam pwm_ctrl_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam pwm_ctrl_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_ctrl_ibuf_1_preio (
            .PADOEN(N__4874),
            .PADOUT(N__4873),
            .PADIN(N__4872),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_ctrl_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_prescale_ibuf_2_iopad (
            .OE(N__4865),
            .DIN(N__4864),
            .DOUT(N__4863),
            .PACKAGEPIN(pwm_prescale[2]));
    defparam pwm_prescale_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam pwm_prescale_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_prescale_ibuf_2_preio (
            .PADOEN(N__4865),
            .PADOUT(N__4864),
            .PADIN(N__4863),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_prescale_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_10_iopad (
            .OE(N__4856),
            .DIN(N__4855),
            .DOUT(N__4854),
            .PACKAGEPIN(pwm_lout[10]));
    defparam pwm_lout_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_10_preio (
            .PADOEN(N__4856),
            .PADOUT(N__4855),
            .PADIN(N__4854),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_8_iopad (
            .OE(N__4847),
            .DIN(N__4846),
            .DOUT(N__4845),
            .PACKAGEPIN(pwm_lout[8]));
    defparam pwm_lout_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_8_preio (
            .PADOEN(N__4847),
            .PADOUT(N__4846),
            .PADIN(N__4845),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_10_iopad (
            .OE(N__4838),
            .DIN(N__4837),
            .DOUT(N__4836),
            .PACKAGEPIN(pwm_hout[10]));
    defparam pwm_hout_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_10_preio (
            .PADOEN(N__4838),
            .PADOUT(N__4837),
            .PADIN(N__4836),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_6_iopad (
            .OE(N__4829),
            .DIN(N__4828),
            .DOUT(N__4827),
            .PACKAGEPIN(pwm_hout[6]));
    defparam pwm_hout_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_6_preio (
            .PADOEN(N__4829),
            .PADOUT(N__4828),
            .PADIN(N__4827),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_0_iopad (
            .OE(N__4820),
            .DIN(N__4819),
            .DOUT(N__4818),
            .PACKAGEPIN(pwm_lout[0]));
    defparam pwm_lout_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_0_preio (
            .PADOEN(N__4820),
            .PADOUT(N__4819),
            .PADIN(N__4818),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_3_iopad (
            .OE(N__4811),
            .DIN(N__4810),
            .DOUT(N__4809),
            .PACKAGEPIN(pwm_hout[3]));
    defparam pwm_hout_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_3_preio (
            .PADOEN(N__4811),
            .PADOUT(N__4810),
            .PADIN(N__4809),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_5_iopad (
            .OE(N__4802),
            .DIN(N__4801),
            .DOUT(N__4800),
            .PACKAGEPIN(pwm_lout[5]));
    defparam pwm_lout_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_5_preio (
            .PADOEN(N__4802),
            .PADOUT(N__4801),
            .PADIN(N__4800),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_8_iopad (
            .OE(N__4793),
            .DIN(N__4792),
            .DOUT(N__4791),
            .PACKAGEPIN(pwm_hout[8]));
    defparam pwm_hout_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_8_preio (
            .PADOEN(N__4793),
            .PADOUT(N__4792),
            .PADIN(N__4791),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_prescale_ibuf_0_iopad (
            .OE(N__4784),
            .DIN(N__4783),
            .DOUT(N__4782),
            .PACKAGEPIN(pwm_prescale[0]));
    defparam pwm_prescale_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam pwm_prescale_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_prescale_ibuf_0_preio (
            .PADOEN(N__4784),
            .PADOUT(N__4783),
            .PADIN(N__4782),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_prescale_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_hout_ibuf_0_iopad (
            .OE(N__4775),
            .DIN(N__4774),
            .DOUT(N__4773),
            .PACKAGEPIN(pwm_hout[0]));
    defparam pwm_hout_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam pwm_hout_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_hout_ibuf_0_preio (
            .PADOEN(N__4775),
            .PADOUT(N__4774),
            .PADIN(N__4773),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_hout_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_2_iopad (
            .OE(N__4766),
            .DIN(N__4765),
            .DOUT(N__4764),
            .PACKAGEPIN(pwm_lout[2]));
    defparam pwm_lout_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_2_preio (
            .PADOEN(N__4766),
            .PADOUT(N__4765),
            .PADIN(N__4764),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_11_iopad (
            .OE(N__4757),
            .DIN(N__4756),
            .DOUT(N__4755),
            .PACKAGEPIN(pwm_lout[11]));
    defparam pwm_lout_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_11_preio (
            .PADOEN(N__4757),
            .PADOUT(N__4756),
            .PADIN(N__4755),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD pwm_lout_ibuf_7_iopad (
            .OE(N__4748),
            .DIN(N__4747),
            .DOUT(N__4746),
            .PACKAGEPIN(pwm_lout[7]));
    defparam pwm_lout_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam pwm_lout_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO pwm_lout_ibuf_7_preio (
            .PADOEN(N__4748),
            .PADOUT(N__4747),
            .PADIN(N__4746),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(pwm_lout_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1020 (
            .O(N__4729),
            .I(N__4723));
    InMux I__1019 (
            .O(N__4728),
            .I(N__4723));
    LocalMux I__1018 (
            .O(N__4723),
            .I(prescale_stop_p1Z0Z_4));
    InMux I__1017 (
            .O(N__4720),
            .I(N__4717));
    LocalMux I__1016 (
            .O(N__4717),
            .I(N__4713));
    InMux I__1015 (
            .O(N__4716),
            .I(N__4710));
    Odrv4 I__1014 (
            .O(N__4713),
            .I(prescale_cntZ0Z_4));
    LocalMux I__1013 (
            .O(N__4710),
            .I(prescale_cntZ0Z_4));
    InMux I__1012 (
            .O(N__4705),
            .I(N__4702));
    LocalMux I__1011 (
            .O(N__4702),
            .I(prescale_cnt_p1Z0Z_4));
    InMux I__1010 (
            .O(N__4699),
            .I(N__4693));
    InMux I__1009 (
            .O(N__4698),
            .I(N__4690));
    InMux I__1008 (
            .O(N__4697),
            .I(N__4684));
    InMux I__1007 (
            .O(N__4696),
            .I(N__4681));
    LocalMux I__1006 (
            .O(N__4693),
            .I(N__4673));
    LocalMux I__1005 (
            .O(N__4690),
            .I(N__4673));
    InMux I__1004 (
            .O(N__4689),
            .I(N__4668));
    InMux I__1003 (
            .O(N__4688),
            .I(N__4668));
    InMux I__1002 (
            .O(N__4687),
            .I(N__4662));
    LocalMux I__1001 (
            .O(N__4684),
            .I(N__4657));
    LocalMux I__1000 (
            .O(N__4681),
            .I(N__4657));
    InMux I__999 (
            .O(N__4680),
            .I(N__4654));
    InMux I__998 (
            .O(N__4679),
            .I(N__4649));
    InMux I__997 (
            .O(N__4678),
            .I(N__4649));
    Span4Mux_v I__996 (
            .O(N__4673),
            .I(N__4643));
    LocalMux I__995 (
            .O(N__4668),
            .I(N__4643));
    InMux I__994 (
            .O(N__4667),
            .I(N__4636));
    InMux I__993 (
            .O(N__4666),
            .I(N__4636));
    InMux I__992 (
            .O(N__4665),
            .I(N__4636));
    LocalMux I__991 (
            .O(N__4662),
            .I(N__4629));
    Span4Mux_v I__990 (
            .O(N__4657),
            .I(N__4629));
    LocalMux I__989 (
            .O(N__4654),
            .I(N__4629));
    LocalMux I__988 (
            .O(N__4649),
            .I(N__4626));
    InMux I__987 (
            .O(N__4648),
            .I(N__4623));
    Span4Mux_h I__986 (
            .O(N__4643),
            .I(N__4620));
    LocalMux I__985 (
            .O(N__4636),
            .I(N__4615));
    Span4Mux_h I__984 (
            .O(N__4629),
            .I(N__4615));
    Span12Mux_h I__983 (
            .O(N__4626),
            .I(N__4610));
    LocalMux I__982 (
            .O(N__4623),
            .I(N__4610));
    Odrv4 I__981 (
            .O(N__4620),
            .I(pwm_prescale_p1Z0Z_2));
    Odrv4 I__980 (
            .O(N__4615),
            .I(pwm_prescale_p1Z0Z_2));
    Odrv12 I__979 (
            .O(N__4610),
            .I(pwm_prescale_p1Z0Z_2));
    CascadeMux I__978 (
            .O(N__4603),
            .I(N__4600));
    InMux I__977 (
            .O(N__4600),
            .I(N__4588));
    InMux I__976 (
            .O(N__4599),
            .I(N__4588));
    InMux I__975 (
            .O(N__4598),
            .I(N__4585));
    InMux I__974 (
            .O(N__4597),
            .I(N__4582));
    InMux I__973 (
            .O(N__4596),
            .I(N__4579));
    InMux I__972 (
            .O(N__4595),
            .I(N__4576));
    InMux I__971 (
            .O(N__4594),
            .I(N__4569));
    InMux I__970 (
            .O(N__4593),
            .I(N__4566));
    LocalMux I__969 (
            .O(N__4588),
            .I(N__4563));
    LocalMux I__968 (
            .O(N__4585),
            .I(N__4556));
    LocalMux I__967 (
            .O(N__4582),
            .I(N__4556));
    LocalMux I__966 (
            .O(N__4579),
            .I(N__4556));
    LocalMux I__965 (
            .O(N__4576),
            .I(N__4553));
    InMux I__964 (
            .O(N__4575),
            .I(N__4550));
    InMux I__963 (
            .O(N__4574),
            .I(N__4545));
    InMux I__962 (
            .O(N__4573),
            .I(N__4545));
    InMux I__961 (
            .O(N__4572),
            .I(N__4542));
    LocalMux I__960 (
            .O(N__4569),
            .I(N__4537));
    LocalMux I__959 (
            .O(N__4566),
            .I(N__4537));
    Span4Mux_v I__958 (
            .O(N__4563),
            .I(N__4532));
    Span4Mux_v I__957 (
            .O(N__4556),
            .I(N__4532));
    Odrv12 I__956 (
            .O(N__4553),
            .I(pwm_prescale_p1Z0Z_1));
    LocalMux I__955 (
            .O(N__4550),
            .I(pwm_prescale_p1Z0Z_1));
    LocalMux I__954 (
            .O(N__4545),
            .I(pwm_prescale_p1Z0Z_1));
    LocalMux I__953 (
            .O(N__4542),
            .I(pwm_prescale_p1Z0Z_1));
    Odrv4 I__952 (
            .O(N__4537),
            .I(pwm_prescale_p1Z0Z_1));
    Odrv4 I__951 (
            .O(N__4532),
            .I(pwm_prescale_p1Z0Z_1));
    InMux I__950 (
            .O(N__4519),
            .I(N__4516));
    LocalMux I__949 (
            .O(N__4516),
            .I(N__4513));
    Odrv4 I__948 (
            .O(N__4513),
            .I(prescale_cnt_p1Z0Z_13));
    InMux I__947 (
            .O(N__4510),
            .I(N__4507));
    LocalMux I__946 (
            .O(N__4507),
            .I(prescale_cnt_p1Z0Z_12));
    InMux I__945 (
            .O(N__4504),
            .I(N__4501));
    LocalMux I__944 (
            .O(N__4501),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_26));
    InMux I__943 (
            .O(N__4498),
            .I(N__4495));
    LocalMux I__942 (
            .O(N__4495),
            .I(prescale_stop_1_8));
    InMux I__941 (
            .O(N__4492),
            .I(N__4481));
    InMux I__940 (
            .O(N__4491),
            .I(N__4481));
    InMux I__939 (
            .O(N__4490),
            .I(N__4481));
    InMux I__938 (
            .O(N__4489),
            .I(N__4475));
    InMux I__937 (
            .O(N__4488),
            .I(N__4472));
    LocalMux I__936 (
            .O(N__4481),
            .I(N__4469));
    InMux I__935 (
            .O(N__4480),
            .I(N__4466));
    InMux I__934 (
            .O(N__4479),
            .I(N__4463));
    InMux I__933 (
            .O(N__4478),
            .I(N__4458));
    LocalMux I__932 (
            .O(N__4475),
            .I(N__4453));
    LocalMux I__931 (
            .O(N__4472),
            .I(N__4453));
    Span4Mux_v I__930 (
            .O(N__4469),
            .I(N__4450));
    LocalMux I__929 (
            .O(N__4466),
            .I(N__4445));
    LocalMux I__928 (
            .O(N__4463),
            .I(N__4445));
    InMux I__927 (
            .O(N__4462),
            .I(N__4440));
    InMux I__926 (
            .O(N__4461),
            .I(N__4440));
    LocalMux I__925 (
            .O(N__4458),
            .I(N__4435));
    Span4Mux_v I__924 (
            .O(N__4453),
            .I(N__4435));
    Span4Mux_v I__923 (
            .O(N__4450),
            .I(N__4427));
    Span4Mux_h I__922 (
            .O(N__4445),
            .I(N__4427));
    LocalMux I__921 (
            .O(N__4440),
            .I(N__4427));
    Span4Mux_h I__920 (
            .O(N__4435),
            .I(N__4424));
    InMux I__919 (
            .O(N__4434),
            .I(N__4421));
    Odrv4 I__918 (
            .O(N__4427),
            .I(pwm_prescale_p1Z0Z_0));
    Odrv4 I__917 (
            .O(N__4424),
            .I(pwm_prescale_p1Z0Z_0));
    LocalMux I__916 (
            .O(N__4421),
            .I(pwm_prescale_p1Z0Z_0));
    InMux I__915 (
            .O(N__4414),
            .I(N__4411));
    LocalMux I__914 (
            .O(N__4411),
            .I(prescale_stop_p1Z0Z_13));
    ClkMux I__913 (
            .O(N__4408),
            .I(N__4333));
    ClkMux I__912 (
            .O(N__4407),
            .I(N__4333));
    ClkMux I__911 (
            .O(N__4406),
            .I(N__4333));
    ClkMux I__910 (
            .O(N__4405),
            .I(N__4333));
    ClkMux I__909 (
            .O(N__4404),
            .I(N__4333));
    ClkMux I__908 (
            .O(N__4403),
            .I(N__4333));
    ClkMux I__907 (
            .O(N__4402),
            .I(N__4333));
    ClkMux I__906 (
            .O(N__4401),
            .I(N__4333));
    ClkMux I__905 (
            .O(N__4400),
            .I(N__4333));
    ClkMux I__904 (
            .O(N__4399),
            .I(N__4333));
    ClkMux I__903 (
            .O(N__4398),
            .I(N__4333));
    ClkMux I__902 (
            .O(N__4397),
            .I(N__4333));
    ClkMux I__901 (
            .O(N__4396),
            .I(N__4333));
    ClkMux I__900 (
            .O(N__4395),
            .I(N__4333));
    ClkMux I__899 (
            .O(N__4394),
            .I(N__4333));
    ClkMux I__898 (
            .O(N__4393),
            .I(N__4333));
    ClkMux I__897 (
            .O(N__4392),
            .I(N__4333));
    ClkMux I__896 (
            .O(N__4391),
            .I(N__4333));
    ClkMux I__895 (
            .O(N__4390),
            .I(N__4333));
    ClkMux I__894 (
            .O(N__4389),
            .I(N__4333));
    ClkMux I__893 (
            .O(N__4388),
            .I(N__4333));
    ClkMux I__892 (
            .O(N__4387),
            .I(N__4333));
    ClkMux I__891 (
            .O(N__4386),
            .I(N__4333));
    ClkMux I__890 (
            .O(N__4385),
            .I(N__4333));
    ClkMux I__889 (
            .O(N__4384),
            .I(N__4333));
    GlobalMux I__888 (
            .O(N__4333),
            .I(N__4330));
    gio2CtrlBuf I__887 (
            .O(N__4330),
            .I(clk_c_g));
    SRMux I__886 (
            .O(N__4327),
            .I(N__4252));
    SRMux I__885 (
            .O(N__4326),
            .I(N__4252));
    SRMux I__884 (
            .O(N__4325),
            .I(N__4252));
    SRMux I__883 (
            .O(N__4324),
            .I(N__4252));
    SRMux I__882 (
            .O(N__4323),
            .I(N__4252));
    SRMux I__881 (
            .O(N__4322),
            .I(N__4252));
    SRMux I__880 (
            .O(N__4321),
            .I(N__4252));
    SRMux I__879 (
            .O(N__4320),
            .I(N__4252));
    SRMux I__878 (
            .O(N__4319),
            .I(N__4252));
    SRMux I__877 (
            .O(N__4318),
            .I(N__4252));
    SRMux I__876 (
            .O(N__4317),
            .I(N__4252));
    SRMux I__875 (
            .O(N__4316),
            .I(N__4252));
    SRMux I__874 (
            .O(N__4315),
            .I(N__4252));
    SRMux I__873 (
            .O(N__4314),
            .I(N__4252));
    SRMux I__872 (
            .O(N__4313),
            .I(N__4252));
    SRMux I__871 (
            .O(N__4312),
            .I(N__4252));
    SRMux I__870 (
            .O(N__4311),
            .I(N__4252));
    SRMux I__869 (
            .O(N__4310),
            .I(N__4252));
    SRMux I__868 (
            .O(N__4309),
            .I(N__4252));
    SRMux I__867 (
            .O(N__4308),
            .I(N__4252));
    SRMux I__866 (
            .O(N__4307),
            .I(N__4252));
    SRMux I__865 (
            .O(N__4306),
            .I(N__4252));
    SRMux I__864 (
            .O(N__4305),
            .I(N__4252));
    SRMux I__863 (
            .O(N__4304),
            .I(N__4252));
    SRMux I__862 (
            .O(N__4303),
            .I(N__4252));
    GlobalMux I__861 (
            .O(N__4252),
            .I(N__4249));
    gio2CtrlBuf I__860 (
            .O(N__4249),
            .I(reset_c_g));
    InMux I__859 (
            .O(N__4246),
            .I(N__4243));
    LocalMux I__858 (
            .O(N__4243),
            .I(N__4240));
    Odrv12 I__857 (
            .O(N__4240),
            .I(prescale_cnt_p1Z0Z_5));
    InMux I__856 (
            .O(N__4237),
            .I(N__4234));
    LocalMux I__855 (
            .O(N__4234),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_6));
    InMux I__854 (
            .O(N__4231),
            .I(N__4228));
    LocalMux I__853 (
            .O(N__4228),
            .I(N__4224));
    InMux I__852 (
            .O(N__4227),
            .I(N__4221));
    Odrv12 I__851 (
            .O(N__4224),
            .I(prescale_stop_p1Z0Z_14));
    LocalMux I__850 (
            .O(N__4221),
            .I(prescale_stop_p1Z0Z_14));
    InMux I__849 (
            .O(N__4216),
            .I(N__4213));
    LocalMux I__848 (
            .O(N__4213),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_36));
    InMux I__847 (
            .O(N__4210),
            .I(N__4207));
    LocalMux I__846 (
            .O(N__4207),
            .I(N__4204));
    Span4Mux_v I__845 (
            .O(N__4204),
            .I(N__4200));
    InMux I__844 (
            .O(N__4203),
            .I(N__4197));
    Odrv4 I__843 (
            .O(N__4200),
            .I(prescale_cntZ0Z_12));
    LocalMux I__842 (
            .O(N__4197),
            .I(prescale_cntZ0Z_12));
    InMux I__841 (
            .O(N__4192),
            .I(N__4189));
    LocalMux I__840 (
            .O(N__4189),
            .I(N__4185));
    InMux I__839 (
            .O(N__4188),
            .I(N__4182));
    Odrv4 I__838 (
            .O(N__4185),
            .I(prescale_cntZ0Z_16));
    LocalMux I__837 (
            .O(N__4182),
            .I(prescale_cntZ0Z_16));
    InMux I__836 (
            .O(N__4177),
            .I(N__4174));
    LocalMux I__835 (
            .O(N__4174),
            .I(prescale_cnt_p1Z0Z_16));
    CascadeMux I__834 (
            .O(N__4171),
            .I(N__4168));
    InMux I__833 (
            .O(N__4168),
            .I(N__4165));
    LocalMux I__832 (
            .O(N__4165),
            .I(prescale_stop_p1Z0Z_5));
    InMux I__831 (
            .O(N__4162),
            .I(N__4159));
    LocalMux I__830 (
            .O(N__4159),
            .I(prescale_stop_1_7));
    InMux I__829 (
            .O(N__4156),
            .I(N__4153));
    LocalMux I__828 (
            .O(N__4153),
            .I(N__4150));
    Span4Mux_h I__827 (
            .O(N__4150),
            .I(N__4146));
    InMux I__826 (
            .O(N__4149),
            .I(N__4143));
    Odrv4 I__825 (
            .O(N__4146),
            .I(prescale_cntZ0Z_3));
    LocalMux I__824 (
            .O(N__4143),
            .I(prescale_cntZ0Z_3));
    InMux I__823 (
            .O(N__4138),
            .I(N__4135));
    LocalMux I__822 (
            .O(N__4135),
            .I(prescale_cnt_p1Z0Z_3));
    InMux I__821 (
            .O(N__4132),
            .I(N__4129));
    LocalMux I__820 (
            .O(N__4129),
            .I(N__4126));
    Span4Mux_h I__819 (
            .O(N__4126),
            .I(N__4122));
    InMux I__818 (
            .O(N__4125),
            .I(N__4119));
    Odrv4 I__817 (
            .O(N__4122),
            .I(prescale_cntZ0Z_2));
    LocalMux I__816 (
            .O(N__4119),
            .I(prescale_cntZ0Z_2));
    InMux I__815 (
            .O(N__4114),
            .I(N__4111));
    LocalMux I__814 (
            .O(N__4111),
            .I(prescale_cnt_p1Z0Z_2));
    InMux I__813 (
            .O(N__4108),
            .I(N__4105));
    LocalMux I__812 (
            .O(N__4105),
            .I(N__4102));
    Span4Mux_h I__811 (
            .O(N__4102),
            .I(N__4098));
    InMux I__810 (
            .O(N__4101),
            .I(N__4095));
    Odrv4 I__809 (
            .O(N__4098),
            .I(prescale_cntZ0Z_13));
    LocalMux I__808 (
            .O(N__4095),
            .I(prescale_cntZ0Z_13));
    InMux I__807 (
            .O(N__4090),
            .I(N__4087));
    LocalMux I__806 (
            .O(N__4087),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_1));
    InMux I__805 (
            .O(N__4084),
            .I(N__4081));
    LocalMux I__804 (
            .O(N__4081),
            .I(N__4078));
    Span4Mux_v I__803 (
            .O(N__4078),
            .I(N__4075));
    Odrv4 I__802 (
            .O(N__4075),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_11));
    InMux I__801 (
            .O(N__4072),
            .I(N__4069));
    LocalMux I__800 (
            .O(N__4069),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_16));
    InMux I__799 (
            .O(N__4066),
            .I(N__4063));
    LocalMux I__798 (
            .O(N__4063),
            .I(N__4060));
    Span4Mux_v I__797 (
            .O(N__4060),
            .I(N__4057));
    Odrv4 I__796 (
            .O(N__4057),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_21));
    InMux I__795 (
            .O(N__4054),
            .I(N__4051));
    LocalMux I__794 (
            .O(N__4051),
            .I(N__4048));
    Odrv12 I__793 (
            .O(N__4048),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_31));
    InMux I__792 (
            .O(N__4045),
            .I(proc_pwm_cnt_prescale_cnt10));
    InMux I__791 (
            .O(N__4042),
            .I(N__4036));
    InMux I__790 (
            .O(N__4041),
            .I(N__4036));
    LocalMux I__789 (
            .O(N__4036),
            .I(N__4033));
    Odrv12 I__788 (
            .O(N__4033),
            .I(proc_pwm_cnt_prescale_cnt10_THRU_CO));
    InMux I__787 (
            .O(N__4030),
            .I(N__4027));
    LocalMux I__786 (
            .O(N__4027),
            .I(N__4024));
    Odrv12 I__785 (
            .O(N__4024),
            .I(pwm_prescale_c_1));
    InMux I__784 (
            .O(N__4021),
            .I(N__4018));
    LocalMux I__783 (
            .O(N__4018),
            .I(N__4015));
    Span4Mux_v I__782 (
            .O(N__4015),
            .I(N__4012));
    Span4Mux_h I__781 (
            .O(N__4012),
            .I(N__4009));
    Sp12to4 I__780 (
            .O(N__4009),
            .I(N__4006));
    Odrv12 I__779 (
            .O(N__4006),
            .I(pwm_lout_c_5));
    InMux I__778 (
            .O(N__4003),
            .I(N__4000));
    LocalMux I__777 (
            .O(N__4000),
            .I(N__3997));
    Odrv12 I__776 (
            .O(N__3997),
            .I(pwm_lout_p1Z0Z_5));
    CascadeMux I__775 (
            .O(N__3994),
            .I(N__3991));
    InMux I__774 (
            .O(N__3991),
            .I(N__3988));
    LocalMux I__773 (
            .O(N__3988),
            .I(prescale_stop_p1Z0Z_8));
    InMux I__772 (
            .O(N__3985),
            .I(N__3982));
    LocalMux I__771 (
            .O(N__3982),
            .I(N__3979));
    Span4Mux_h I__770 (
            .O(N__3979),
            .I(N__3975));
    InMux I__769 (
            .O(N__3978),
            .I(N__3972));
    Odrv4 I__768 (
            .O(N__3975),
            .I(prescale_cntZ0Z_8));
    LocalMux I__767 (
            .O(N__3972),
            .I(prescale_cntZ0Z_8));
    InMux I__766 (
            .O(N__3967),
            .I(N__3964));
    LocalMux I__765 (
            .O(N__3964),
            .I(prescale_cnt_p1Z0Z_8));
    InMux I__764 (
            .O(N__3961),
            .I(N__3958));
    LocalMux I__763 (
            .O(N__3958),
            .I(N__3955));
    Span4Mux_h I__762 (
            .O(N__3955),
            .I(N__3951));
    InMux I__761 (
            .O(N__3954),
            .I(N__3948));
    Odrv4 I__760 (
            .O(N__3951),
            .I(prescale_cntZ0Z_9));
    LocalMux I__759 (
            .O(N__3948),
            .I(prescale_cntZ0Z_9));
    InMux I__758 (
            .O(N__3943),
            .I(N__3940));
    LocalMux I__757 (
            .O(N__3940),
            .I(prescale_cnt_p1Z0Z_9));
    InMux I__756 (
            .O(N__3937),
            .I(N__3931));
    InMux I__755 (
            .O(N__3936),
            .I(N__3931));
    LocalMux I__754 (
            .O(N__3931),
            .I(prescale_stop_p1Z0Z_2));
    CascadeMux I__753 (
            .O(N__3928),
            .I(N__3925));
    InMux I__752 (
            .O(N__3925),
            .I(N__3922));
    LocalMux I__751 (
            .O(N__3922),
            .I(prescale_stop_p1Z0Z_3));
    InMux I__750 (
            .O(N__3919),
            .I(N__3916));
    LocalMux I__749 (
            .O(N__3916),
            .I(N__3913));
    Span4Mux_h I__748 (
            .O(N__3913),
            .I(N__3910));
    Odrv4 I__747 (
            .O(N__3910),
            .I(proc_pwm_cnt_prescale_cnt10_0_N_41));
    CascadeMux I__746 (
            .O(N__3907),
            .I(N__3904));
    InMux I__745 (
            .O(N__3904),
            .I(N__3901));
    LocalMux I__744 (
            .O(N__3901),
            .I(prescale_stop_p1Z0Z_1));
    InMux I__743 (
            .O(N__3898),
            .I(N__3895));
    LocalMux I__742 (
            .O(N__3895),
            .I(N__3892));
    Span4Mux_h I__741 (
            .O(N__3892),
            .I(N__3889));
    Span4Mux_v I__740 (
            .O(N__3889),
            .I(N__3886));
    Span4Mux_v I__739 (
            .O(N__3886),
            .I(N__3883));
    Odrv4 I__738 (
            .O(N__3883),
            .I(pwm_lout_c_4));
    InMux I__737 (
            .O(N__3880),
            .I(N__3877));
    LocalMux I__736 (
            .O(N__3877),
            .I(N__3874));
    Odrv12 I__735 (
            .O(N__3874),
            .I(pwm_lout_p1Z0Z_4));
    InMux I__734 (
            .O(N__3871),
            .I(N__3868));
    LocalMux I__733 (
            .O(N__3868),
            .I(N__3865));
    Span4Mux_v I__732 (
            .O(N__3865),
            .I(N__3861));
    InMux I__731 (
            .O(N__3864),
            .I(N__3858));
    Odrv4 I__730 (
            .O(N__3861),
            .I(prescale_cntZ0Z_5));
    LocalMux I__729 (
            .O(N__3858),
            .I(prescale_cntZ0Z_5));
    CascadeMux I__728 (
            .O(N__3853),
            .I(N__3850));
    InMux I__727 (
            .O(N__3850),
            .I(N__3847));
    LocalMux I__726 (
            .O(N__3847),
            .I(prescale_stop_p1Z0Z_15));
    InMux I__725 (
            .O(N__3844),
            .I(N__3841));
    LocalMux I__724 (
            .O(N__3841),
            .I(N__3838));
    Span12Mux_v I__723 (
            .O(N__3838),
            .I(N__3834));
    InMux I__722 (
            .O(N__3837),
            .I(N__3831));
    Odrv12 I__721 (
            .O(N__3834),
            .I(prescale_cntZ0Z_14));
    LocalMux I__720 (
            .O(N__3831),
            .I(prescale_cntZ0Z_14));
    InMux I__719 (
            .O(N__3826),
            .I(N__3823));
    LocalMux I__718 (
            .O(N__3823),
            .I(prescale_cnt_p1Z0Z_14));
    InMux I__717 (
            .O(N__3820),
            .I(N__3817));
    LocalMux I__716 (
            .O(N__3817),
            .I(N__3814));
    Span4Mux_h I__715 (
            .O(N__3814),
            .I(N__3811));
    Span4Mux_v I__714 (
            .O(N__3811),
            .I(N__3807));
    InMux I__713 (
            .O(N__3810),
            .I(N__3804));
    Odrv4 I__712 (
            .O(N__3807),
            .I(prescale_cntZ0Z_15));
    LocalMux I__711 (
            .O(N__3804),
            .I(prescale_cntZ0Z_15));
    InMux I__710 (
            .O(N__3799),
            .I(N__3796));
    LocalMux I__709 (
            .O(N__3796),
            .I(prescale_cnt_p1Z0Z_15));
    InMux I__708 (
            .O(N__3793),
            .I(prescale_cnt_cry_8));
    InMux I__707 (
            .O(N__3790),
            .I(N__3787));
    LocalMux I__706 (
            .O(N__3787),
            .I(N__3783));
    InMux I__705 (
            .O(N__3786),
            .I(N__3780));
    Odrv12 I__704 (
            .O(N__3783),
            .I(prescale_cntZ0Z_10));
    LocalMux I__703 (
            .O(N__3780),
            .I(prescale_cntZ0Z_10));
    InMux I__702 (
            .O(N__3775),
            .I(prescale_cnt_cry_9));
    InMux I__701 (
            .O(N__3772),
            .I(N__3769));
    LocalMux I__700 (
            .O(N__3769),
            .I(N__3765));
    InMux I__699 (
            .O(N__3768),
            .I(N__3762));
    Odrv12 I__698 (
            .O(N__3765),
            .I(prescale_cntZ0Z_11));
    LocalMux I__697 (
            .O(N__3762),
            .I(prescale_cntZ0Z_11));
    InMux I__696 (
            .O(N__3757),
            .I(prescale_cnt_cry_10));
    InMux I__695 (
            .O(N__3754),
            .I(prescale_cnt_cry_11));
    InMux I__694 (
            .O(N__3751),
            .I(prescale_cnt_cry_12));
    InMux I__693 (
            .O(N__3748),
            .I(prescale_cnt_cry_13));
    InMux I__692 (
            .O(N__3745),
            .I(prescale_cnt_cry_14));
    InMux I__691 (
            .O(N__3742),
            .I(N__3724));
    InMux I__690 (
            .O(N__3741),
            .I(N__3715));
    InMux I__689 (
            .O(N__3740),
            .I(N__3715));
    InMux I__688 (
            .O(N__3739),
            .I(N__3715));
    InMux I__687 (
            .O(N__3738),
            .I(N__3715));
    InMux I__686 (
            .O(N__3737),
            .I(N__3706));
    InMux I__685 (
            .O(N__3736),
            .I(N__3706));
    InMux I__684 (
            .O(N__3735),
            .I(N__3706));
    InMux I__683 (
            .O(N__3734),
            .I(N__3706));
    InMux I__682 (
            .O(N__3733),
            .I(N__3699));
    InMux I__681 (
            .O(N__3732),
            .I(N__3699));
    InMux I__680 (
            .O(N__3731),
            .I(N__3699));
    InMux I__679 (
            .O(N__3730),
            .I(N__3690));
    InMux I__678 (
            .O(N__3729),
            .I(N__3690));
    InMux I__677 (
            .O(N__3728),
            .I(N__3690));
    InMux I__676 (
            .O(N__3727),
            .I(N__3690));
    LocalMux I__675 (
            .O(N__3724),
            .I(N_8));
    LocalMux I__674 (
            .O(N__3715),
            .I(N_8));
    LocalMux I__673 (
            .O(N__3706),
            .I(N_8));
    LocalMux I__672 (
            .O(N__3699),
            .I(N_8));
    LocalMux I__671 (
            .O(N__3690),
            .I(N_8));
    InMux I__670 (
            .O(N__3679),
            .I(bfn_3_14_0_));
    InMux I__669 (
            .O(N__3676),
            .I(N__3668));
    InMux I__668 (
            .O(N__3675),
            .I(N__3668));
    InMux I__667 (
            .O(N__3674),
            .I(N__3663));
    InMux I__666 (
            .O(N__3673),
            .I(N__3663));
    LocalMux I__665 (
            .O(N__3668),
            .I(prescale_stop_p1Z0Z_0));
    LocalMux I__664 (
            .O(N__3663),
            .I(prescale_stop_p1Z0Z_0));
    InMux I__663 (
            .O(N__3658),
            .I(N__3654));
    InMux I__662 (
            .O(N__3657),
            .I(N__3651));
    LocalMux I__661 (
            .O(N__3654),
            .I(prescale_cntZ0Z_1));
    LocalMux I__660 (
            .O(N__3651),
            .I(prescale_cntZ0Z_1));
    InMux I__659 (
            .O(N__3646),
            .I(prescale_cnt_cry_0));
    InMux I__658 (
            .O(N__3643),
            .I(prescale_cnt_cry_1));
    InMux I__657 (
            .O(N__3640),
            .I(prescale_cnt_cry_2));
    InMux I__656 (
            .O(N__3637),
            .I(prescale_cnt_cry_3));
    InMux I__655 (
            .O(N__3634),
            .I(prescale_cnt_cry_4));
    InMux I__654 (
            .O(N__3631),
            .I(N__3628));
    LocalMux I__653 (
            .O(N__3628),
            .I(N__3624));
    InMux I__652 (
            .O(N__3627),
            .I(N__3621));
    Odrv12 I__651 (
            .O(N__3624),
            .I(prescale_cntZ0Z_6));
    LocalMux I__650 (
            .O(N__3621),
            .I(prescale_cntZ0Z_6));
    InMux I__649 (
            .O(N__3616),
            .I(prescale_cnt_cry_5));
    InMux I__648 (
            .O(N__3613),
            .I(N__3610));
    LocalMux I__647 (
            .O(N__3610),
            .I(N__3606));
    InMux I__646 (
            .O(N__3609),
            .I(N__3603));
    Odrv12 I__645 (
            .O(N__3606),
            .I(prescale_cntZ0Z_7));
    LocalMux I__644 (
            .O(N__3603),
            .I(prescale_cntZ0Z_7));
    InMux I__643 (
            .O(N__3598),
            .I(prescale_cnt_cry_6));
    InMux I__642 (
            .O(N__3595),
            .I(bfn_3_13_0_));
    InMux I__641 (
            .O(N__3592),
            .I(N__3588));
    InMux I__640 (
            .O(N__3591),
            .I(N__3585));
    LocalMux I__639 (
            .O(N__3588),
            .I(N__3580));
    LocalMux I__638 (
            .O(N__3585),
            .I(N__3580));
    Odrv4 I__637 (
            .O(N__3580),
            .I(pwm_ctrl_p1Z0Z_0));
    InMux I__636 (
            .O(N__3577),
            .I(N__3573));
    InMux I__635 (
            .O(N__3576),
            .I(N__3570));
    LocalMux I__634 (
            .O(N__3573),
            .I(N__3567));
    LocalMux I__633 (
            .O(N__3570),
            .I(N__3564));
    Odrv4 I__632 (
            .O(N__3567),
            .I(pwm_ctrl_p1Z0Z_1));
    Odrv4 I__631 (
            .O(N__3564),
            .I(pwm_ctrl_p1Z0Z_1));
    CascadeMux I__630 (
            .O(N__3559),
            .I(pwm_loc_1_sqmuxa_cascade_));
    CascadeMux I__629 (
            .O(N__3556),
            .I(un1_pwm_loc8_1_0_cascade_));
    CEMux I__628 (
            .O(N__3553),
            .I(N__3549));
    CEMux I__627 (
            .O(N__3552),
            .I(N__3546));
    LocalMux I__626 (
            .O(N__3549),
            .I(pwm_cnte_0_i));
    LocalMux I__625 (
            .O(N__3546),
            .I(pwm_cnte_0_i));
    InMux I__624 (
            .O(N__3541),
            .I(N__3538));
    LocalMux I__623 (
            .O(N__3538),
            .I(un1_pwm_loc8_1_0));
    CascadeMux I__622 (
            .O(N__3535),
            .I(N__3531));
    CascadeMux I__621 (
            .O(N__3534),
            .I(N__3526));
    InMux I__620 (
            .O(N__3531),
            .I(N__3519));
    InMux I__619 (
            .O(N__3530),
            .I(N__3519));
    InMux I__618 (
            .O(N__3529),
            .I(N__3519));
    InMux I__617 (
            .O(N__3526),
            .I(N__3516));
    LocalMux I__616 (
            .O(N__3519),
            .I(N__3513));
    LocalMux I__615 (
            .O(N__3516),
            .I(N__3510));
    Odrv4 I__614 (
            .O(N__3513),
            .I(prescale_tickZ0));
    Odrv4 I__613 (
            .O(N__3510),
            .I(prescale_tickZ0));
    InMux I__612 (
            .O(N__3505),
            .I(N__3502));
    LocalMux I__611 (
            .O(N__3502),
            .I(pwm_loc_1_sqmuxa));
    InMux I__610 (
            .O(N__3499),
            .I(N__3496));
    LocalMux I__609 (
            .O(N__3496),
            .I(pwm_loc_0_sqmuxa_1));
    CascadeMux I__608 (
            .O(N__3493),
            .I(pwm_loc_1_sqmuxa_1_cascade_));
    InMux I__607 (
            .O(N__3490),
            .I(N__3487));
    LocalMux I__606 (
            .O(N__3487),
            .I(N__3484));
    Span4Mux_h I__605 (
            .O(N__3484),
            .I(N__3481));
    Span4Mux_v I__604 (
            .O(N__3481),
            .I(N__3477));
    InMux I__603 (
            .O(N__3480),
            .I(N__3474));
    Odrv4 I__602 (
            .O(N__3477),
            .I(pwm_locZ0));
    LocalMux I__601 (
            .O(N__3474),
            .I(pwm_locZ0));
    InMux I__600 (
            .O(N__3469),
            .I(N__3464));
    InMux I__599 (
            .O(N__3468),
            .I(N__3459));
    InMux I__598 (
            .O(N__3467),
            .I(N__3459));
    LocalMux I__597 (
            .O(N__3464),
            .I(proc_pwm_fsm_pwm_loc20_THRU_CO));
    LocalMux I__596 (
            .O(N__3459),
            .I(proc_pwm_fsm_pwm_loc20_THRU_CO));
    InMux I__595 (
            .O(N__3454),
            .I(N__3451));
    LocalMux I__594 (
            .O(N__3451),
            .I(N_87));
    CascadeMux I__593 (
            .O(N__3448),
            .I(N__3445));
    InMux I__592 (
            .O(N__3445),
            .I(N__3437));
    InMux I__591 (
            .O(N__3444),
            .I(N__3434));
    InMux I__590 (
            .O(N__3443),
            .I(N__3425));
    InMux I__589 (
            .O(N__3442),
            .I(N__3425));
    InMux I__588 (
            .O(N__3441),
            .I(N__3425));
    InMux I__587 (
            .O(N__3440),
            .I(N__3425));
    LocalMux I__586 (
            .O(N__3437),
            .I(pwm_toglZ0));
    LocalMux I__585 (
            .O(N__3434),
            .I(pwm_toglZ0));
    LocalMux I__584 (
            .O(N__3425),
            .I(pwm_toglZ0));
    InMux I__583 (
            .O(N__3418),
            .I(N__3406));
    InMux I__582 (
            .O(N__3417),
            .I(N__3406));
    InMux I__581 (
            .O(N__3416),
            .I(N__3406));
    InMux I__580 (
            .O(N__3415),
            .I(N__3406));
    LocalMux I__579 (
            .O(N__3406),
            .I(N__3403));
    Odrv4 I__578 (
            .O(N__3403),
            .I(N_86));
    CascadeMux I__577 (
            .O(N__3400),
            .I(N_87_cascade_));
    InMux I__576 (
            .O(N__3397),
            .I(N__3388));
    InMux I__575 (
            .O(N__3396),
            .I(N__3388));
    InMux I__574 (
            .O(N__3395),
            .I(N__3388));
    LocalMux I__573 (
            .O(N__3388),
            .I(N__3384));
    InMux I__572 (
            .O(N__3387),
            .I(N__3381));
    Span4Mux_h I__571 (
            .O(N__3384),
            .I(N__3378));
    LocalMux I__570 (
            .O(N__3381),
            .I(proc_pwm_fsm_pwm_loc8_THRU_CO));
    Odrv4 I__569 (
            .O(N__3378),
            .I(proc_pwm_fsm_pwm_loc8_THRU_CO));
    InMux I__568 (
            .O(N__3373),
            .I(N__3359));
    InMux I__567 (
            .O(N__3372),
            .I(N__3359));
    InMux I__566 (
            .O(N__3371),
            .I(N__3359));
    InMux I__565 (
            .O(N__3370),
            .I(N__3359));
    InMux I__564 (
            .O(N__3369),
            .I(N__3348));
    InMux I__563 (
            .O(N__3368),
            .I(N__3348));
    LocalMux I__562 (
            .O(N__3359),
            .I(N__3345));
    InMux I__561 (
            .O(N__3358),
            .I(N__3340));
    InMux I__560 (
            .O(N__3357),
            .I(N__3340));
    InMux I__559 (
            .O(N__3356),
            .I(N__3331));
    InMux I__558 (
            .O(N__3355),
            .I(N__3331));
    InMux I__557 (
            .O(N__3354),
            .I(N__3331));
    InMux I__556 (
            .O(N__3353),
            .I(N__3331));
    LocalMux I__555 (
            .O(N__3348),
            .I(N_78_0_i));
    Odrv4 I__554 (
            .O(N__3345),
            .I(N_78_0_i));
    LocalMux I__553 (
            .O(N__3340),
            .I(N_78_0_i));
    LocalMux I__552 (
            .O(N__3331),
            .I(N_78_0_i));
    InMux I__551 (
            .O(N__3322),
            .I(N__3318));
    InMux I__550 (
            .O(N__3321),
            .I(N__3315));
    LocalMux I__549 (
            .O(N__3318),
            .I(prescale_cntZ0Z_0));
    LocalMux I__548 (
            .O(N__3315),
            .I(prescale_cntZ0Z_0));
    InMux I__547 (
            .O(N__3310),
            .I(N__3307));
    LocalMux I__546 (
            .O(N__3307),
            .I(prescale_cnt_s_0));
    InMux I__545 (
            .O(N__3304),
            .I(bfn_3_12_0_));
    InMux I__544 (
            .O(N__3301),
            .I(N__3298));
    LocalMux I__543 (
            .O(N__3298),
            .I(prescale_stop_p1Z0Z_6));
    InMux I__542 (
            .O(N__3295),
            .I(N__3292));
    LocalMux I__541 (
            .O(N__3292),
            .I(prescale_cnt_p1Z0Z_7));
    CascadeMux I__540 (
            .O(N__3289),
            .I(N__3286));
    InMux I__539 (
            .O(N__3286),
            .I(N__3283));
    LocalMux I__538 (
            .O(N__3283),
            .I(prescale_stop_p1Z0Z_7));
    InMux I__537 (
            .O(N__3280),
            .I(N__3277));
    LocalMux I__536 (
            .O(N__3277),
            .I(prescale_cnt_p1Z0Z_6));
    InMux I__535 (
            .O(N__3274),
            .I(N__3271));
    LocalMux I__534 (
            .O(N__3271),
            .I(prescale_stop_p1Z0Z_10));
    InMux I__533 (
            .O(N__3268),
            .I(N__3265));
    LocalMux I__532 (
            .O(N__3265),
            .I(prescale_cnt_p1Z0Z_11));
    InMux I__531 (
            .O(N__3262),
            .I(N__3259));
    LocalMux I__530 (
            .O(N__3259),
            .I(prescale_cnt_p1Z0Z_10));
    InMux I__529 (
            .O(N__3256),
            .I(N__3251));
    InMux I__528 (
            .O(N__3255),
            .I(N__3248));
    InMux I__527 (
            .O(N__3254),
            .I(N__3245));
    LocalMux I__526 (
            .O(N__3251),
            .I(pwm_cntZ0Z_1));
    LocalMux I__525 (
            .O(N__3248),
            .I(pwm_cntZ0Z_1));
    LocalMux I__524 (
            .O(N__3245),
            .I(pwm_cntZ0Z_1));
    InMux I__523 (
            .O(N__3238),
            .I(N__3235));
    LocalMux I__522 (
            .O(N__3235),
            .I(N__3232));
    Odrv4 I__521 (
            .O(N__3232),
            .I(pwm_lout_p1Z0Z_1));
    CascadeMux I__520 (
            .O(N__3229),
            .I(N__3225));
    InMux I__519 (
            .O(N__3228),
            .I(N__3221));
    InMux I__518 (
            .O(N__3225),
            .I(N__3218));
    InMux I__517 (
            .O(N__3224),
            .I(N__3215));
    LocalMux I__516 (
            .O(N__3221),
            .I(pwm_cntZ0Z_0));
    LocalMux I__515 (
            .O(N__3218),
            .I(pwm_cntZ0Z_0));
    LocalMux I__514 (
            .O(N__3215),
            .I(pwm_cntZ0Z_0));
    InMux I__513 (
            .O(N__3208),
            .I(N__3205));
    LocalMux I__512 (
            .O(N__3205),
            .I(pwm_lout_p1Z0Z_0));
    CascadeMux I__511 (
            .O(N__3202),
            .I(N__3199));
    InMux I__510 (
            .O(N__3199),
            .I(N__3196));
    LocalMux I__509 (
            .O(N__3196),
            .I(proc_pwm_fsm_pwm_loc20_0_N_26));
    CascadeMux I__508 (
            .O(N__3193),
            .I(N__3189));
    InMux I__507 (
            .O(N__3192),
            .I(N__3185));
    InMux I__506 (
            .O(N__3189),
            .I(N__3182));
    InMux I__505 (
            .O(N__3188),
            .I(N__3179));
    LocalMux I__504 (
            .O(N__3185),
            .I(pwm_cntZ0Z_5));
    LocalMux I__503 (
            .O(N__3182),
            .I(pwm_cntZ0Z_5));
    LocalMux I__502 (
            .O(N__3179),
            .I(pwm_cntZ0Z_5));
    InMux I__501 (
            .O(N__3172),
            .I(N__3167));
    InMux I__500 (
            .O(N__3171),
            .I(N__3164));
    InMux I__499 (
            .O(N__3170),
            .I(N__3161));
    LocalMux I__498 (
            .O(N__3167),
            .I(pwm_cntZ0Z_4));
    LocalMux I__497 (
            .O(N__3164),
            .I(pwm_cntZ0Z_4));
    LocalMux I__496 (
            .O(N__3161),
            .I(pwm_cntZ0Z_4));
    CascadeMux I__495 (
            .O(N__3154),
            .I(N__3151));
    InMux I__494 (
            .O(N__3151),
            .I(N__3148));
    LocalMux I__493 (
            .O(N__3148),
            .I(proc_pwm_fsm_pwm_loc20_0_N_16));
    InMux I__492 (
            .O(N__3145),
            .I(N__3142));
    LocalMux I__491 (
            .O(N__3142),
            .I(N__3139));
    Span4Mux_h I__490 (
            .O(N__3139),
            .I(N__3136));
    Span4Mux_v I__489 (
            .O(N__3136),
            .I(N__3133));
    Span4Mux_v I__488 (
            .O(N__3133),
            .I(N__3130));
    Odrv4 I__487 (
            .O(N__3130),
            .I(pwm_lout_c_11));
    CascadeMux I__486 (
            .O(N__3127),
            .I(N__3124));
    InMux I__485 (
            .O(N__3124),
            .I(N__3121));
    LocalMux I__484 (
            .O(N__3121),
            .I(pwm_lout_p1Z0Z_11));
    InMux I__483 (
            .O(N__3118),
            .I(N__3115));
    LocalMux I__482 (
            .O(N__3115),
            .I(N__3112));
    Span12Mux_v I__481 (
            .O(N__3112),
            .I(N__3109));
    Odrv12 I__480 (
            .O(N__3109),
            .I(pwm_lout_c_10));
    InMux I__479 (
            .O(N__3106),
            .I(N__3103));
    LocalMux I__478 (
            .O(N__3103),
            .I(pwm_lout_p1Z0Z_10));
    InMux I__477 (
            .O(N__3100),
            .I(N__3097));
    LocalMux I__476 (
            .O(N__3097),
            .I(N__3094));
    Sp12to4 I__475 (
            .O(N__3094),
            .I(N__3091));
    Span12Mux_v I__474 (
            .O(N__3091),
            .I(N__3088));
    Odrv12 I__473 (
            .O(N__3088),
            .I(pwm_lout_c_1));
    InMux I__472 (
            .O(N__3085),
            .I(N__3082));
    LocalMux I__471 (
            .O(N__3082),
            .I(N__3079));
    Span4Mux_v I__470 (
            .O(N__3079),
            .I(N__3076));
    Sp12to4 I__469 (
            .O(N__3076),
            .I(N__3073));
    Odrv12 I__468 (
            .O(N__3073),
            .I(pwm_ctrl_c_1));
    InMux I__467 (
            .O(N__3070),
            .I(N__3067));
    LocalMux I__466 (
            .O(N__3067),
            .I(N__3064));
    Span12Mux_h I__465 (
            .O(N__3064),
            .I(N__3061));
    Span12Mux_v I__464 (
            .O(N__3061),
            .I(N__3058));
    Odrv12 I__463 (
            .O(N__3058),
            .I(pwm_lout_c_0));
    InMux I__462 (
            .O(N__3055),
            .I(pwm_cnt_cry_9));
    InMux I__461 (
            .O(N__3052),
            .I(pwm_cnt_cry_10));
    CascadeMux I__460 (
            .O(N__3049),
            .I(N_8_cascade_));
    InMux I__459 (
            .O(N__3046),
            .I(N__3043));
    LocalMux I__458 (
            .O(N__3043),
            .I(prescale_cnt_p1Z0Z_0));
    InMux I__457 (
            .O(N__3040),
            .I(N__3037));
    LocalMux I__456 (
            .O(N__3037),
            .I(prescale_cnt_p1Z0Z_1));
    InMux I__455 (
            .O(N__3034),
            .I(N__3025));
    InMux I__454 (
            .O(N__3033),
            .I(N__3025));
    InMux I__453 (
            .O(N__3032),
            .I(N__3025));
    LocalMux I__452 (
            .O(N__3025),
            .I(N_38));
    InMux I__451 (
            .O(N__3022),
            .I(N__3017));
    InMux I__450 (
            .O(N__3021),
            .I(N__3014));
    InMux I__449 (
            .O(N__3020),
            .I(N__3011));
    LocalMux I__448 (
            .O(N__3017),
            .I(N__3008));
    LocalMux I__447 (
            .O(N__3014),
            .I(pwm_cntZ0Z_11));
    LocalMux I__446 (
            .O(N__3011),
            .I(pwm_cntZ0Z_11));
    Odrv4 I__445 (
            .O(N__3008),
            .I(pwm_cntZ0Z_11));
    InMux I__444 (
            .O(N__3001),
            .I(N__2996));
    InMux I__443 (
            .O(N__3000),
            .I(N__2993));
    InMux I__442 (
            .O(N__2999),
            .I(N__2990));
    LocalMux I__441 (
            .O(N__2996),
            .I(N__2987));
    LocalMux I__440 (
            .O(N__2993),
            .I(pwm_cntZ0Z_10));
    LocalMux I__439 (
            .O(N__2990),
            .I(pwm_cntZ0Z_10));
    Odrv4 I__438 (
            .O(N__2987),
            .I(pwm_cntZ0Z_10));
    CascadeMux I__437 (
            .O(N__2980),
            .I(N__2977));
    InMux I__436 (
            .O(N__2977),
            .I(N__2974));
    LocalMux I__435 (
            .O(N__2974),
            .I(N__2971));
    Odrv12 I__434 (
            .O(N__2971),
            .I(proc_pwm_fsm_pwm_loc20_0_N_1));
    InMux I__433 (
            .O(N__2968),
            .I(N__2963));
    InMux I__432 (
            .O(N__2967),
            .I(N__2960));
    InMux I__431 (
            .O(N__2966),
            .I(N__2957));
    LocalMux I__430 (
            .O(N__2963),
            .I(pwm_cntZ0Z_2));
    LocalMux I__429 (
            .O(N__2960),
            .I(pwm_cntZ0Z_2));
    LocalMux I__428 (
            .O(N__2957),
            .I(pwm_cntZ0Z_2));
    InMux I__427 (
            .O(N__2950),
            .I(pwm_cnt_cry_1));
    InMux I__426 (
            .O(N__2947),
            .I(N__2942));
    InMux I__425 (
            .O(N__2946),
            .I(N__2937));
    InMux I__424 (
            .O(N__2945),
            .I(N__2937));
    LocalMux I__423 (
            .O(N__2942),
            .I(pwm_cntZ0Z_3));
    LocalMux I__422 (
            .O(N__2937),
            .I(pwm_cntZ0Z_3));
    InMux I__421 (
            .O(N__2932),
            .I(pwm_cnt_cry_2));
    InMux I__420 (
            .O(N__2929),
            .I(pwm_cnt_cry_3));
    InMux I__419 (
            .O(N__2926),
            .I(pwm_cnt_cry_4));
    InMux I__418 (
            .O(N__2923),
            .I(N__2918));
    InMux I__417 (
            .O(N__2922),
            .I(N__2915));
    InMux I__416 (
            .O(N__2921),
            .I(N__2912));
    LocalMux I__415 (
            .O(N__2918),
            .I(pwm_cntZ0Z_6));
    LocalMux I__414 (
            .O(N__2915),
            .I(pwm_cntZ0Z_6));
    LocalMux I__413 (
            .O(N__2912),
            .I(pwm_cntZ0Z_6));
    InMux I__412 (
            .O(N__2905),
            .I(pwm_cnt_cry_5));
    InMux I__411 (
            .O(N__2902),
            .I(N__2897));
    InMux I__410 (
            .O(N__2901),
            .I(N__2894));
    InMux I__409 (
            .O(N__2900),
            .I(N__2891));
    LocalMux I__408 (
            .O(N__2897),
            .I(pwm_cntZ0Z_7));
    LocalMux I__407 (
            .O(N__2894),
            .I(pwm_cntZ0Z_7));
    LocalMux I__406 (
            .O(N__2891),
            .I(pwm_cntZ0Z_7));
    InMux I__405 (
            .O(N__2884),
            .I(pwm_cnt_cry_6));
    InMux I__404 (
            .O(N__2881),
            .I(N__2876));
    InMux I__403 (
            .O(N__2880),
            .I(N__2873));
    InMux I__402 (
            .O(N__2879),
            .I(N__2870));
    LocalMux I__401 (
            .O(N__2876),
            .I(N__2867));
    LocalMux I__400 (
            .O(N__2873),
            .I(pwm_cntZ0Z_8));
    LocalMux I__399 (
            .O(N__2870),
            .I(pwm_cntZ0Z_8));
    Odrv4 I__398 (
            .O(N__2867),
            .I(pwm_cntZ0Z_8));
    InMux I__397 (
            .O(N__2860),
            .I(bfn_2_12_0_));
    InMux I__396 (
            .O(N__2857),
            .I(N__2852));
    InMux I__395 (
            .O(N__2856),
            .I(N__2849));
    InMux I__394 (
            .O(N__2855),
            .I(N__2846));
    LocalMux I__393 (
            .O(N__2852),
            .I(N__2843));
    LocalMux I__392 (
            .O(N__2849),
            .I(pwm_cntZ0Z_9));
    LocalMux I__391 (
            .O(N__2846),
            .I(pwm_cntZ0Z_9));
    Odrv4 I__390 (
            .O(N__2843),
            .I(pwm_cntZ0Z_9));
    InMux I__389 (
            .O(N__2836),
            .I(pwm_cnt_cry_8));
    CascadeMux I__388 (
            .O(N__2833),
            .I(N__2830));
    InMux I__387 (
            .O(N__2830),
            .I(N__2827));
    LocalMux I__386 (
            .O(N__2827),
            .I(proc_pwm_fsm_pwm_loc20_0_N_21));
    CascadeMux I__385 (
            .O(N__2824),
            .I(N__2821));
    InMux I__384 (
            .O(N__2821),
            .I(N__2818));
    LocalMux I__383 (
            .O(N__2818),
            .I(proc_pwm_fsm_pwm_loc20_0_N_6));
    CascadeMux I__382 (
            .O(N__2815),
            .I(N__2812));
    InMux I__381 (
            .O(N__2812),
            .I(N__2809));
    LocalMux I__380 (
            .O(N__2809),
            .I(proc_pwm_fsm_pwm_loc20_0_N_11));
    InMux I__379 (
            .O(N__2806),
            .I(proc_pwm_fsm_pwm_loc20));
    InMux I__378 (
            .O(N__2803),
            .I(bfn_2_11_0_));
    InMux I__377 (
            .O(N__2800),
            .I(pwm_cnt_cry_0));
    InMux I__376 (
            .O(N__2797),
            .I(N__2794));
    LocalMux I__375 (
            .O(N__2794),
            .I(N__2791));
    Span4Mux_v I__374 (
            .O(N__2791),
            .I(N__2788));
    Span4Mux_v I__373 (
            .O(N__2788),
            .I(N__2785));
    Span4Mux_h I__372 (
            .O(N__2785),
            .I(N__2782));
    Odrv4 I__371 (
            .O(N__2782),
            .I(pwm_hout_c_7));
    CascadeMux I__370 (
            .O(N__2779),
            .I(N__2776));
    InMux I__369 (
            .O(N__2776),
            .I(N__2773));
    LocalMux I__368 (
            .O(N__2773),
            .I(N__2770));
    Span4Mux_h I__367 (
            .O(N__2770),
            .I(N__2767));
    Odrv4 I__366 (
            .O(N__2767),
            .I(pwm_hout_p1Z0Z_7));
    InMux I__365 (
            .O(N__2764),
            .I(N__2761));
    LocalMux I__364 (
            .O(N__2761),
            .I(N__2758));
    Span4Mux_h I__363 (
            .O(N__2758),
            .I(N__2755));
    Span4Mux_v I__362 (
            .O(N__2755),
            .I(N__2752));
    Span4Mux_v I__361 (
            .O(N__2752),
            .I(N__2749));
    Odrv4 I__360 (
            .O(N__2749),
            .I(pwm_hout_c_11));
    CascadeMux I__359 (
            .O(N__2746),
            .I(N__2743));
    InMux I__358 (
            .O(N__2743),
            .I(N__2740));
    LocalMux I__357 (
            .O(N__2740),
            .I(pwm_hout_p1Z0Z_11));
    InMux I__356 (
            .O(N__2737),
            .I(N__2734));
    LocalMux I__355 (
            .O(N__2734),
            .I(N__2731));
    Span4Mux_v I__354 (
            .O(N__2731),
            .I(N__2728));
    Span4Mux_h I__353 (
            .O(N__2728),
            .I(N__2725));
    Odrv4 I__352 (
            .O(N__2725),
            .I(pwm_prescale_c_0));
    InMux I__351 (
            .O(N__2722),
            .I(N__2719));
    LocalMux I__350 (
            .O(N__2719),
            .I(N__2716));
    Span4Mux_v I__349 (
            .O(N__2716),
            .I(N__2713));
    Sp12to4 I__348 (
            .O(N__2713),
            .I(N__2710));
    Odrv12 I__347 (
            .O(N__2710),
            .I(pwm_lout_c_7));
    InMux I__346 (
            .O(N__2707),
            .I(N__2704));
    LocalMux I__345 (
            .O(N__2704),
            .I(N__2701));
    Odrv12 I__344 (
            .O(N__2701),
            .I(pwm_lout_p1Z0Z_7));
    InMux I__343 (
            .O(N__2698),
            .I(N__2695));
    LocalMux I__342 (
            .O(N__2695),
            .I(N__2692));
    Span12Mux_v I__341 (
            .O(N__2692),
            .I(N__2689));
    Odrv12 I__340 (
            .O(N__2689),
            .I(pwm_prescale_c_2));
    InMux I__339 (
            .O(N__2686),
            .I(N__2683));
    LocalMux I__338 (
            .O(N__2683),
            .I(N__2680));
    Span12Mux_v I__337 (
            .O(N__2680),
            .I(N__2677));
    Odrv12 I__336 (
            .O(N__2677),
            .I(pwm_lout_c_8));
    InMux I__335 (
            .O(N__2674),
            .I(N__2671));
    LocalMux I__334 (
            .O(N__2671),
            .I(N__2668));
    Span12Mux_v I__333 (
            .O(N__2668),
            .I(N__2665));
    Odrv12 I__332 (
            .O(N__2665),
            .I(pwm_ctrl_c_0));
    CascadeMux I__331 (
            .O(N__2662),
            .I(N__2659));
    InMux I__330 (
            .O(N__2659),
            .I(N__2656));
    LocalMux I__329 (
            .O(N__2656),
            .I(pwm_lout_p1Z0Z_8));
    InMux I__328 (
            .O(N__2653),
            .I(N__2650));
    LocalMux I__327 (
            .O(N__2650),
            .I(pwm_lout_p1Z0Z_9));
    InMux I__326 (
            .O(N__2647),
            .I(N__2644));
    LocalMux I__325 (
            .O(N__2644),
            .I(N__2641));
    Span4Mux_h I__324 (
            .O(N__2641),
            .I(N__2638));
    Span4Mux_v I__323 (
            .O(N__2638),
            .I(N__2635));
    Odrv4 I__322 (
            .O(N__2635),
            .I(pwm_hout_c_0));
    InMux I__321 (
            .O(N__2632),
            .I(N__2629));
    LocalMux I__320 (
            .O(N__2629),
            .I(pwm_hout_p1Z0Z_0));
    InMux I__319 (
            .O(N__2626),
            .I(N__2623));
    LocalMux I__318 (
            .O(N__2623),
            .I(N__2620));
    Span4Mux_v I__317 (
            .O(N__2620),
            .I(N__2617));
    Span4Mux_h I__316 (
            .O(N__2617),
            .I(N__2614));
    Odrv4 I__315 (
            .O(N__2614),
            .I(pwm_hout_c_3));
    CascadeMux I__314 (
            .O(N__2611),
            .I(N__2608));
    InMux I__313 (
            .O(N__2608),
            .I(N__2605));
    LocalMux I__312 (
            .O(N__2605),
            .I(pwm_hout_p1Z0Z_3));
    InMux I__311 (
            .O(N__2602),
            .I(N__2599));
    LocalMux I__310 (
            .O(N__2599),
            .I(N__2596));
    Span12Mux_h I__309 (
            .O(N__2596),
            .I(N__2593));
    Span12Mux_v I__308 (
            .O(N__2593),
            .I(N__2590));
    Odrv12 I__307 (
            .O(N__2590),
            .I(pwm_lout_c_2));
    CascadeMux I__306 (
            .O(N__2587),
            .I(N__2584));
    InMux I__305 (
            .O(N__2584),
            .I(N__2581));
    LocalMux I__304 (
            .O(N__2581),
            .I(pwm_lout_p1Z0Z_2));
    InMux I__303 (
            .O(N__2578),
            .I(N__2575));
    LocalMux I__302 (
            .O(N__2575),
            .I(N__2572));
    Span4Mux_h I__301 (
            .O(N__2572),
            .I(N__2569));
    Span4Mux_v I__300 (
            .O(N__2569),
            .I(N__2566));
    Odrv4 I__299 (
            .O(N__2566),
            .I(pwm_hout_c_1));
    CascadeMux I__298 (
            .O(N__2563),
            .I(N__2560));
    InMux I__297 (
            .O(N__2560),
            .I(N__2557));
    LocalMux I__296 (
            .O(N__2557),
            .I(pwm_hout_p1Z0Z_1));
    InMux I__295 (
            .O(N__2554),
            .I(N__2551));
    LocalMux I__294 (
            .O(N__2551),
            .I(N__2548));
    Span4Mux_v I__293 (
            .O(N__2548),
            .I(N__2545));
    Span4Mux_v I__292 (
            .O(N__2545),
            .I(N__2542));
    Span4Mux_h I__291 (
            .O(N__2542),
            .I(N__2539));
    Odrv4 I__290 (
            .O(N__2539),
            .I(pwm_hout_c_2));
    InMux I__289 (
            .O(N__2536),
            .I(N__2533));
    LocalMux I__288 (
            .O(N__2533),
            .I(pwm_hout_p1Z0Z_2));
    InMux I__287 (
            .O(N__2530),
            .I(N__2527));
    LocalMux I__286 (
            .O(N__2527),
            .I(N__2524));
    Odrv12 I__285 (
            .O(N__2524),
            .I(pwm_lout_c_3));
    InMux I__284 (
            .O(N__2521),
            .I(N__2518));
    LocalMux I__283 (
            .O(N__2518),
            .I(pwm_lout_p1Z0Z_3));
    InMux I__282 (
            .O(N__2515),
            .I(N__2512));
    LocalMux I__281 (
            .O(N__2512),
            .I(N__2509));
    Odrv12 I__280 (
            .O(N__2509),
            .I(proc_pwm_fsm_pwm_loc8_0_N_1));
    InMux I__279 (
            .O(N__2506),
            .I(N__2503));
    LocalMux I__278 (
            .O(N__2503),
            .I(N__2500));
    Sp12to4 I__277 (
            .O(N__2500),
            .I(N__2497));
    Span12Mux_v I__276 (
            .O(N__2497),
            .I(N__2494));
    Odrv12 I__275 (
            .O(N__2494),
            .I(pwm_hout_c_6));
    InMux I__274 (
            .O(N__2491),
            .I(N__2488));
    LocalMux I__273 (
            .O(N__2488),
            .I(N__2485));
    Odrv4 I__272 (
            .O(N__2485),
            .I(pwm_hout_p1Z0Z_6));
    InMux I__271 (
            .O(N__2482),
            .I(N__2479));
    LocalMux I__270 (
            .O(N__2479),
            .I(N__2476));
    Span4Mux_v I__269 (
            .O(N__2476),
            .I(N__2473));
    Span4Mux_v I__268 (
            .O(N__2473),
            .I(N__2470));
    Span4Mux_h I__267 (
            .O(N__2470),
            .I(N__2467));
    Odrv4 I__266 (
            .O(N__2467),
            .I(pwm_hout_c_10));
    InMux I__265 (
            .O(N__2464),
            .I(N__2461));
    LocalMux I__264 (
            .O(N__2461),
            .I(pwm_hout_p1Z0Z_10));
    CascadeMux I__263 (
            .O(N__2458),
            .I(N__2455));
    InMux I__262 (
            .O(N__2455),
            .I(N__2452));
    LocalMux I__261 (
            .O(N__2452),
            .I(pwm_lout_p1Z0Z_6));
    CascadeMux I__260 (
            .O(N__2449),
            .I(N__2446));
    InMux I__259 (
            .O(N__2446),
            .I(N__2443));
    LocalMux I__258 (
            .O(N__2443),
            .I(proc_pwm_fsm_pwm_loc8_0_N_26));
    InMux I__257 (
            .O(N__2440),
            .I(N__2437));
    LocalMux I__256 (
            .O(N__2437),
            .I(proc_pwm_fsm_pwm_loc8_0_N_6));
    InMux I__255 (
            .O(N__2434),
            .I(N__2431));
    LocalMux I__254 (
            .O(N__2431),
            .I(proc_pwm_fsm_pwm_loc8_0_N_16));
    InMux I__253 (
            .O(N__2428),
            .I(N__2425));
    LocalMux I__252 (
            .O(N__2425),
            .I(proc_pwm_fsm_pwm_loc8_0_N_21));
    InMux I__251 (
            .O(N__2422),
            .I(N__2419));
    LocalMux I__250 (
            .O(N__2419),
            .I(N__2416));
    Odrv4 I__249 (
            .O(N__2416),
            .I(pwm_hout_p1Z0Z_8));
    CascadeMux I__248 (
            .O(N__2413),
            .I(N__2410));
    InMux I__247 (
            .O(N__2410),
            .I(N__2407));
    LocalMux I__246 (
            .O(N__2407),
            .I(N__2404));
    Span4Mux_v I__245 (
            .O(N__2404),
            .I(N__2401));
    Odrv4 I__244 (
            .O(N__2401),
            .I(pwm_hout_p1Z0Z_9));
    InMux I__243 (
            .O(N__2398),
            .I(N__2395));
    LocalMux I__242 (
            .O(N__2395),
            .I(proc_pwm_fsm_pwm_loc8_0_N_11));
    InMux I__241 (
            .O(N__2392),
            .I(N__2389));
    LocalMux I__240 (
            .O(N__2389),
            .I(N__2386));
    Span4Mux_v I__239 (
            .O(N__2386),
            .I(N__2383));
    Sp12to4 I__238 (
            .O(N__2383),
            .I(N__2380));
    Span12Mux_h I__237 (
            .O(N__2380),
            .I(N__2377));
    Odrv12 I__236 (
            .O(N__2377),
            .I(pwm_hout_c_5));
    CascadeMux I__235 (
            .O(N__2374),
            .I(N__2371));
    InMux I__234 (
            .O(N__2371),
            .I(N__2368));
    LocalMux I__233 (
            .O(N__2368),
            .I(pwm_hout_p1Z0Z_5));
    InMux I__232 (
            .O(N__2365),
            .I(N__2362));
    LocalMux I__231 (
            .O(N__2362),
            .I(N__2359));
    Span4Mux_h I__230 (
            .O(N__2359),
            .I(N__2356));
    Span4Mux_v I__229 (
            .O(N__2356),
            .I(N__2353));
    Span4Mux_v I__228 (
            .O(N__2353),
            .I(N__2350));
    Span4Mux_v I__227 (
            .O(N__2350),
            .I(N__2347));
    Odrv4 I__226 (
            .O(N__2347),
            .I(pwm_hout_c_4));
    InMux I__225 (
            .O(N__2344),
            .I(N__2341));
    LocalMux I__224 (
            .O(N__2341),
            .I(pwm_hout_p1Z0Z_4));
    InMux I__223 (
            .O(N__2338),
            .I(N__2335));
    LocalMux I__222 (
            .O(N__2335),
            .I(N__2332));
    Sp12to4 I__221 (
            .O(N__2332),
            .I(N__2329));
    Span12Mux_v I__220 (
            .O(N__2329),
            .I(N__2326));
    Odrv12 I__219 (
            .O(N__2326),
            .I(pwm_hout_c_9));
    InMux I__218 (
            .O(N__2323),
            .I(N__2320));
    LocalMux I__217 (
            .O(N__2320),
            .I(N__2317));
    Span4Mux_v I__216 (
            .O(N__2317),
            .I(N__2314));
    Span4Mux_v I__215 (
            .O(N__2314),
            .I(N__2311));
    Span4Mux_v I__214 (
            .O(N__2311),
            .I(N__2308));
    Sp12to4 I__213 (
            .O(N__2308),
            .I(N__2305));
    Odrv12 I__212 (
            .O(N__2305),
            .I(pwm_hout_c_8));
    InMux I__211 (
            .O(N__2302),
            .I(proc_pwm_fsm_pwm_loc8));
    IoInMux I__210 (
            .O(N__2299),
            .I(N__2296));
    LocalMux I__209 (
            .O(N__2296),
            .I(N__2293));
    IoSpan4Mux I__208 (
            .O(N__2293),
            .I(N__2290));
    Span4Mux_s3_h I__207 (
            .O(N__2290),
            .I(N__2287));
    Odrv4 I__206 (
            .O(N__2287),
            .I(pwm_pin_c));
    InMux I__205 (
            .O(N__2284),
            .I(N__2281));
    LocalMux I__204 (
            .O(N__2281),
            .I(N__2278));
    Span4Mux_v I__203 (
            .O(N__2278),
            .I(N__2275));
    Span4Mux_v I__202 (
            .O(N__2275),
            .I(N__2272));
    Sp12to4 I__201 (
            .O(N__2272),
            .I(N__2269));
    Odrv12 I__200 (
            .O(N__2269),
            .I(pwm_lout_c_9));
    InMux I__199 (
            .O(N__2266),
            .I(N__2263));
    LocalMux I__198 (
            .O(N__2263),
            .I(N__2260));
    Span4Mux_h I__197 (
            .O(N__2260),
            .I(N__2257));
    Sp12to4 I__196 (
            .O(N__2257),
            .I(N__2254));
    Span12Mux_v I__195 (
            .O(N__2254),
            .I(N__2251));
    Odrv12 I__194 (
            .O(N__2251),
            .I(pwm_lout_c_6));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_5_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_12_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_7),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_12_0_ (
            .carryinitin(pwm_cnt_cry_7),
            .carryinitout(bfn_2_12_0_));
    defparam IN_MUX_bfv_3_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_12_0_));
    defparam IN_MUX_bfv_3_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_13_0_ (
            .carryinitin(prescale_cnt_cry_7),
            .carryinitout(bfn_3_13_0_));
    defparam IN_MUX_bfv_3_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_14_0_ (
            .carryinitin(prescale_cnt_cry_15),
            .carryinitout(bfn_3_14_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam pwm_pinZ0_LC_1_6_6.C_ON=1'b0;
    defparam pwm_pinZ0_LC_1_6_6.SEQ_MODE=4'b1010;
    defparam pwm_pinZ0_LC_1_6_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_pinZ0_LC_1_6_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3490),
            .lcout(pwm_pin_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4393),
            .ce(),
            .sr(N__4317));
    defparam pwm_lout_p1_9_LC_1_8_0.C_ON=1'b0;
    defparam pwm_lout_p1_9_LC_1_8_0.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_9_LC_1_8_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_lout_p1_9_LC_1_8_0 (
            .in0(N__2284),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_lout_p1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4385),
            .ce(),
            .sr(N__4308));
    defparam pwm_lout_p1_6_LC_1_9_0.C_ON=1'b0;
    defparam pwm_lout_p1_6_LC_1_9_0.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_6_LC_1_9_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_lout_p1_6_LC_1_9_0 (
            .in0(N__2266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_lout_p1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4384),
            .ce(),
            .sr(N__4306));
    defparam pwm_hout_p1_9_LC_1_9_2.C_ON=1'b0;
    defparam pwm_hout_p1_9_LC_1_9_2.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_9_LC_1_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_9_LC_1_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2338),
            .lcout(pwm_hout_p1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4384),
            .ce(),
            .sr(N__4306));
    defparam pwm_hout_p1_8_LC_1_9_7.C_ON=1'b0;
    defparam pwm_hout_p1_8_LC_1_9_7.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_8_LC_1_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_8_LC_1_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2323),
            .lcout(pwm_hout_p1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4384),
            .ce(),
            .sr(N__4306));
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_LC_1_10_0.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_LC_1_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_1_c_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(proc_pwm_fsm_pwm_loc8_0_data_tmp_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_LC_1_10_1.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_LC_1_10_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_9_c_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(N__2428),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc8_0_data_tmp_0),
            .carryout(proc_pwm_fsm_pwm_loc8_0_data_tmp_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_LC_1_10_2.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_LC_1_10_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_15_c_LC_1_10_2 (
            .in0(_gnd_net_),
            .in1(N__2434),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc8_0_data_tmp_1),
            .carryout(proc_pwm_fsm_pwm_loc8_0_data_tmp_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_LC_1_10_3.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_LC_1_10_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_LC_1_10_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_27_c_LC_1_10_3 (
            .in0(_gnd_net_),
            .in1(N__2440),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc8_0_data_tmp_2),
            .carryout(proc_pwm_fsm_pwm_loc8_0_data_tmp_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_LC_1_10_4.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_LC_1_10_4.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_LC_1_10_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_21_c_LC_1_10_4 (
            .in0(_gnd_net_),
            .in1(N__2398),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc8_0_data_tmp_3),
            .carryout(proc_pwm_fsm_pwm_loc8_0_data_tmp_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_LC_1_10_5.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_LC_1_10_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_LC_1_10_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_33_c_LC_1_10_5 (
            .in0(_gnd_net_),
            .in1(N__2515),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc8_0_data_tmp_4),
            .carryout(proc_pwm_fsm_pwm_loc8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_THRU_LUT4_0_LC_1_10_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_THRU_LUT4_0_LC_1_10_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_THRU_LUT4_0_LC_1_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_THRU_LUT4_0_LC_1_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2302),
            .lcout(proc_pwm_fsm_pwm_loc8_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_RNO_LC_1_10_7.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_RNO_LC_1_10_7.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_RNO_LC_1_10_7.LUT_INIT=16'b1001000000001001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_27_c_RNO_LC_1_10_7 (
            .in0(N__2707),
            .in1(N__2901),
            .in2(N__2458),
            .in3(N__2921),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_RNO_LC_1_11_0.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_RNO_LC_1_11_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_1_c_RNO_LC_1_11_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_1_c_RNO_LC_1_11_0 (
            .in0(N__2632),
            .in1(N__3254),
            .in2(N__2563),
            .in3(N__3224),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_RNO_LC_1_11_1.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_RNO_LC_1_11_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_27_c_RNO_LC_1_11_1.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_27_c_RNO_LC_1_11_1 (
            .in0(N__2491),
            .in1(N__2900),
            .in2(N__2779),
            .in3(N__2922),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_RNO_LC_1_11_2.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_RNO_LC_1_11_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_RNO_LC_1_11_2.LUT_INIT=16'b1000010000100001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_9_c_RNO_LC_1_11_2 (
            .in0(N__2967),
            .in1(N__2946),
            .in2(N__2587),
            .in3(N__2521),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_RNO_LC_1_11_3.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_RNO_LC_1_11_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_15_c_RNO_LC_1_11_3.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_15_c_RNO_LC_1_11_3 (
            .in0(N__2344),
            .in1(N__3188),
            .in2(N__2374),
            .in3(N__3171),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_RNO_LC_1_11_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_RNO_LC_1_11_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_9_c_RNO_LC_1_11_6.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_9_c_RNO_LC_1_11_6 (
            .in0(N__2536),
            .in1(N__2945),
            .in2(N__2611),
            .in3(N__2966),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_RNO_LC_1_11_7.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_RNO_LC_1_11_7.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_21_c_RNO_LC_1_11_7.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_21_c_RNO_LC_1_11_7 (
            .in0(N__2422),
            .in1(N__2855),
            .in2(N__2413),
            .in3(N__2879),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_hout_p1_5_LC_1_12_0.C_ON=1'b0;
    defparam pwm_hout_p1_5_LC_1_12_0.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_5_LC_1_12_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_hout_p1_5_LC_1_12_0 (
            .in0(N__2392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_hout_p1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_hout_p1_4_LC_1_12_1.C_ON=1'b0;
    defparam pwm_hout_p1_4_LC_1_12_1.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_4_LC_1_12_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_hout_p1_4_LC_1_12_1 (
            .in0(N__2365),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_hout_p1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_hout_p1_0_LC_1_12_2.C_ON=1'b0;
    defparam pwm_hout_p1_0_LC_1_12_2.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_0_LC_1_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_0_LC_1_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2647),
            .lcout(pwm_hout_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_hout_p1_3_LC_1_12_3.C_ON=1'b0;
    defparam pwm_hout_p1_3_LC_1_12_3.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_3_LC_1_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_3_LC_1_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2626),
            .lcout(pwm_hout_p1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_lout_p1_2_LC_1_12_4.C_ON=1'b0;
    defparam pwm_lout_p1_2_LC_1_12_4.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_2_LC_1_12_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_lout_p1_2_LC_1_12_4 (
            .in0(N__2602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_lout_p1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_hout_p1_1_LC_1_12_5.C_ON=1'b0;
    defparam pwm_hout_p1_1_LC_1_12_5.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_1_LC_1_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_hout_p1_1_LC_1_12_5 (
            .in0(N__2578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_hout_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_hout_p1_2_LC_1_12_6.C_ON=1'b0;
    defparam pwm_hout_p1_2_LC_1_12_6.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_2_LC_1_12_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_hout_p1_2_LC_1_12_6 (
            .in0(N__2554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_hout_p1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam pwm_lout_p1_3_LC_1_12_7.C_ON=1'b0;
    defparam pwm_lout_p1_3_LC_1_12_7.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_3_LC_1_12_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_lout_p1_3_LC_1_12_7 (
            .in0(N__2530),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_lout_p1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4386),
            .ce(),
            .sr(N__4304));
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNO_LC_1_13_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNO_LC_1_13_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNO_LC_1_13_6.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_33_c_RNO_LC_1_13_6 (
            .in0(N__2464),
            .in1(N__3020),
            .in2(N__2746),
            .in3(N__2999),
            .lcout(proc_pwm_fsm_pwm_loc8_0_N_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_hout_p1_6_LC_1_14_0.C_ON=1'b0;
    defparam pwm_hout_p1_6_LC_1_14_0.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_6_LC_1_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_6_LC_1_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2506),
            .lcout(pwm_hout_p1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_hout_p1_10_LC_1_14_2.C_ON=1'b0;
    defparam pwm_hout_p1_10_LC_1_14_2.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_10_LC_1_14_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_10_LC_1_14_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2482),
            .lcout(pwm_hout_p1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_hout_p1_7_LC_1_14_3.C_ON=1'b0;
    defparam pwm_hout_p1_7_LC_1_14_3.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_7_LC_1_14_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_7_LC_1_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2797),
            .lcout(pwm_hout_p1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_hout_p1_11_LC_1_14_4.C_ON=1'b0;
    defparam pwm_hout_p1_11_LC_1_14_4.SEQ_MODE=4'b1010;
    defparam pwm_hout_p1_11_LC_1_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_hout_p1_11_LC_1_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2764),
            .lcout(pwm_hout_p1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_prescale_p1_0_LC_1_14_6.C_ON=1'b0;
    defparam pwm_prescale_p1_0_LC_1_14_6.SEQ_MODE=4'b1010;
    defparam pwm_prescale_p1_0_LC_1_14_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_prescale_p1_0_LC_1_14_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2737),
            .lcout(pwm_prescale_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_lout_p1_7_LC_1_14_7.C_ON=1'b0;
    defparam pwm_lout_p1_7_LC_1_14_7.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_7_LC_1_14_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_7_LC_1_14_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2722),
            .lcout(pwm_lout_p1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4394),
            .ce(),
            .sr(N__4309));
    defparam pwm_prescale_p1_2_LC_2_7_7.C_ON=1'b0;
    defparam pwm_prescale_p1_2_LC_2_7_7.SEQ_MODE=4'b1010;
    defparam pwm_prescale_p1_2_LC_2_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_prescale_p1_2_LC_2_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2698),
            .lcout(pwm_prescale_p1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4395),
            .ce(),
            .sr(N__4318));
    defparam pwm_lout_p1_8_LC_2_8_2.C_ON=1'b0;
    defparam pwm_lout_p1_8_LC_2_8_2.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_8_LC_2_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_8_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2686),
            .lcout(pwm_lout_p1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4388),
            .ce(),
            .sr(N__4313));
    defparam pwm_ctrl_p1_0_LC_2_8_5.C_ON=1'b0;
    defparam pwm_ctrl_p1_0_LC_2_8_5.SEQ_MODE=4'b1010;
    defparam pwm_ctrl_p1_0_LC_2_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_ctrl_p1_0_LC_2_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2674),
            .lcout(pwm_ctrl_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4388),
            .ce(),
            .sr(N__4313));
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_RNO_LC_2_9_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_RNO_LC_2_9_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_RNO_LC_2_9_6.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_21_c_RNO_LC_2_9_6 (
            .in0(N__2857),
            .in1(N__2881),
            .in2(N__2662),
            .in3(N__2653),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_LC_2_10_0.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_LC_2_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_1_c_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3202),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(proc_pwm_fsm_pwm_loc20_0_data_tmp_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_LC_2_10_1.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_LC_2_10_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_9_c_LC_2_10_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_9_c_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2833),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc20_0_data_tmp_0),
            .carryout(proc_pwm_fsm_pwm_loc20_0_data_tmp_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_LC_2_10_2.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_LC_2_10_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_LC_2_10_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_15_c_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3154),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc20_0_data_tmp_1),
            .carryout(proc_pwm_fsm_pwm_loc20_0_data_tmp_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_LC_2_10_3.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_LC_2_10_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_27_c_LC_2_10_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_27_c_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2824),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc20_0_data_tmp_2),
            .carryout(proc_pwm_fsm_pwm_loc20_0_data_tmp_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_LC_2_10_4.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_LC_2_10_4.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_21_c_LC_2_10_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_21_c_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2815),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc20_0_data_tmp_3),
            .carryout(proc_pwm_fsm_pwm_loc20_0_data_tmp_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_LC_2_10_5.C_ON=1'b1;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_LC_2_10_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_LC_2_10_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_33_c_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2980),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_fsm_pwm_loc20_0_data_tmp_4),
            .carryout(proc_pwm_fsm_pwm_loc20),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_THRU_LUT4_0_LC_2_10_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_THRU_LUT4_0_LC_2_10_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_THRU_LUT4_0_LC_2_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_THRU_LUT4_0_LC_2_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2806),
            .lcout(proc_pwm_fsm_pwm_loc20_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_loc_RNO_0_LC_2_10_7.C_ON=1'b0;
    defparam pwm_loc_RNO_0_LC_2_10_7.SEQ_MODE=4'b0000;
    defparam pwm_loc_RNO_0_LC_2_10_7.LUT_INIT=16'b0010000011100000;
    LogicCell40 pwm_loc_RNO_0_LC_2_10_7 (
            .in0(N__3387),
            .in1(N__3444),
            .in2(N__3534),
            .in3(N__3469),
            .lcout(pwm_loc_0_sqmuxa_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_cnt_0_LC_2_11_0.C_ON=1'b1;
    defparam pwm_cnt_0_LC_2_11_0.SEQ_MODE=4'b1010;
    defparam pwm_cnt_0_LC_2_11_0.LUT_INIT=16'b1011101111101110;
    LogicCell40 pwm_cnt_0_LC_2_11_0 (
            .in0(N__3370),
            .in1(N__3228),
            .in2(_gnd_net_),
            .in3(N__2803),
            .lcout(pwm_cntZ0Z_0),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(pwm_cnt_cry_0),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_1_LC_2_11_1.C_ON=1'b1;
    defparam pwm_cnt_1_LC_2_11_1.SEQ_MODE=4'b1010;
    defparam pwm_cnt_1_LC_2_11_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_1_LC_2_11_1 (
            .in0(N__3353),
            .in1(N__3256),
            .in2(_gnd_net_),
            .in3(N__2800),
            .lcout(pwm_cntZ0Z_1),
            .ltout(),
            .carryin(pwm_cnt_cry_0),
            .carryout(pwm_cnt_cry_1),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_2_LC_2_11_2.C_ON=1'b1;
    defparam pwm_cnt_2_LC_2_11_2.SEQ_MODE=4'b1010;
    defparam pwm_cnt_2_LC_2_11_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_2_LC_2_11_2 (
            .in0(N__3371),
            .in1(N__2968),
            .in2(_gnd_net_),
            .in3(N__2950),
            .lcout(pwm_cntZ0Z_2),
            .ltout(),
            .carryin(pwm_cnt_cry_1),
            .carryout(pwm_cnt_cry_2),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_3_LC_2_11_3.C_ON=1'b1;
    defparam pwm_cnt_3_LC_2_11_3.SEQ_MODE=4'b1010;
    defparam pwm_cnt_3_LC_2_11_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_3_LC_2_11_3 (
            .in0(N__3354),
            .in1(N__2947),
            .in2(_gnd_net_),
            .in3(N__2932),
            .lcout(pwm_cntZ0Z_3),
            .ltout(),
            .carryin(pwm_cnt_cry_2),
            .carryout(pwm_cnt_cry_3),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_4_LC_2_11_4.C_ON=1'b1;
    defparam pwm_cnt_4_LC_2_11_4.SEQ_MODE=4'b1010;
    defparam pwm_cnt_4_LC_2_11_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_4_LC_2_11_4 (
            .in0(N__3372),
            .in1(N__3172),
            .in2(_gnd_net_),
            .in3(N__2929),
            .lcout(pwm_cntZ0Z_4),
            .ltout(),
            .carryin(pwm_cnt_cry_3),
            .carryout(pwm_cnt_cry_4),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_5_LC_2_11_5.C_ON=1'b1;
    defparam pwm_cnt_5_LC_2_11_5.SEQ_MODE=4'b1010;
    defparam pwm_cnt_5_LC_2_11_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_5_LC_2_11_5 (
            .in0(N__3355),
            .in1(N__3192),
            .in2(_gnd_net_),
            .in3(N__2926),
            .lcout(pwm_cntZ0Z_5),
            .ltout(),
            .carryin(pwm_cnt_cry_4),
            .carryout(pwm_cnt_cry_5),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_6_LC_2_11_6.C_ON=1'b1;
    defparam pwm_cnt_6_LC_2_11_6.SEQ_MODE=4'b1010;
    defparam pwm_cnt_6_LC_2_11_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_6_LC_2_11_6 (
            .in0(N__3373),
            .in1(N__2923),
            .in2(_gnd_net_),
            .in3(N__2905),
            .lcout(pwm_cntZ0Z_6),
            .ltout(),
            .carryin(pwm_cnt_cry_5),
            .carryout(pwm_cnt_cry_6),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_7_LC_2_11_7.C_ON=1'b1;
    defparam pwm_cnt_7_LC_2_11_7.SEQ_MODE=4'b1010;
    defparam pwm_cnt_7_LC_2_11_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_7_LC_2_11_7 (
            .in0(N__3356),
            .in1(N__2902),
            .in2(_gnd_net_),
            .in3(N__2884),
            .lcout(pwm_cntZ0Z_7),
            .ltout(),
            .carryin(pwm_cnt_cry_6),
            .carryout(pwm_cnt_cry_7),
            .clk(N__4387),
            .ce(N__3552),
            .sr(N__4303));
    defparam pwm_cnt_8_LC_2_12_0.C_ON=1'b1;
    defparam pwm_cnt_8_LC_2_12_0.SEQ_MODE=4'b1010;
    defparam pwm_cnt_8_LC_2_12_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_8_LC_2_12_0 (
            .in0(N__3369),
            .in1(N__2880),
            .in2(_gnd_net_),
            .in3(N__2860),
            .lcout(pwm_cntZ0Z_8),
            .ltout(),
            .carryin(bfn_2_12_0_),
            .carryout(pwm_cnt_cry_8),
            .clk(N__4389),
            .ce(N__3553),
            .sr(N__4307));
    defparam pwm_cnt_9_LC_2_12_1.C_ON=1'b1;
    defparam pwm_cnt_9_LC_2_12_1.SEQ_MODE=4'b1010;
    defparam pwm_cnt_9_LC_2_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_9_LC_2_12_1 (
            .in0(N__3357),
            .in1(N__2856),
            .in2(_gnd_net_),
            .in3(N__2836),
            .lcout(pwm_cntZ0Z_9),
            .ltout(),
            .carryin(pwm_cnt_cry_8),
            .carryout(pwm_cnt_cry_9),
            .clk(N__4389),
            .ce(N__3553),
            .sr(N__4307));
    defparam pwm_cnt_10_LC_2_12_2.C_ON=1'b1;
    defparam pwm_cnt_10_LC_2_12_2.SEQ_MODE=4'b1010;
    defparam pwm_cnt_10_LC_2_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_10_LC_2_12_2 (
            .in0(N__3368),
            .in1(N__3000),
            .in2(_gnd_net_),
            .in3(N__3055),
            .lcout(pwm_cntZ0Z_10),
            .ltout(),
            .carryin(pwm_cnt_cry_9),
            .carryout(pwm_cnt_cry_10),
            .clk(N__4389),
            .ce(N__3553),
            .sr(N__4307));
    defparam pwm_cnt_11_LC_2_12_3.C_ON=1'b0;
    defparam pwm_cnt_11_LC_2_12_3.SEQ_MODE=4'b1010;
    defparam pwm_cnt_11_LC_2_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 pwm_cnt_11_LC_2_12_3 (
            .in0(N__3358),
            .in1(N__3021),
            .in2(_gnd_net_),
            .in3(N__3052),
            .lcout(pwm_cntZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4389),
            .ce(N__3553),
            .sr(N__4307));
    defparam prescale_tick_LC_2_13_0.C_ON=1'b0;
    defparam prescale_tick_LC_2_13_0.SEQ_MODE=4'b1010;
    defparam prescale_tick_LC_2_13_0.LUT_INIT=16'b1110111011001100;
    LogicCell40 prescale_tick_LC_2_13_0 (
            .in0(N__4042),
            .in1(N__3033),
            .in2(_gnd_net_),
            .in3(N__3675),
            .lcout(prescale_tickZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4396),
            .ce(),
            .sr(N__4310));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNIRR0O1_LC_2_13_1.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNIRR0O1_LC_2_13_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNIRR0O1_LC_2_13_1.LUT_INIT=16'b1111111110111011;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNIRR0O1_LC_2_13_1 (
            .in0(N__3032),
            .in1(N__3674),
            .in2(_gnd_net_),
            .in3(N__4041),
            .lcout(N_8),
            .ltout(N_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_0_LC_2_13_2.C_ON=1'b0;
    defparam prescale_cnt_0_LC_2_13_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_0_LC_2_13_2.LUT_INIT=16'b0011101000001010;
    LogicCell40 prescale_cnt_0_LC_2_13_2 (
            .in0(N__3310),
            .in1(N__3034),
            .in2(N__3049),
            .in3(N__3676),
            .lcout(prescale_cntZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4396),
            .ce(),
            .sr(N__4310));
    defparam prescale_cnt_p1_0_LC_2_13_3.C_ON=1'b0;
    defparam prescale_cnt_p1_0_LC_2_13_3.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_0_LC_2_13_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_0_LC_2_13_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3322),
            .lcout(prescale_cnt_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4396),
            .ce(),
            .sr(N__4310));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_RNO_LC_2_13_4.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_RNO_LC_2_13_4.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_RNO_LC_2_13_4.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_1_c_RNO_LC_2_13_4 (
            .in0(N__3673),
            .in1(N__3040),
            .in2(N__3907),
            .in3(N__3046),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_41),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_p1_1_LC_2_13_5.C_ON=1'b0;
    defparam prescale_cnt_p1_1_LC_2_13_5.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_1_LC_2_13_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_1_LC_2_13_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3658),
            .lcout(prescale_cnt_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4396),
            .ce(),
            .sr(N__4310));
    defparam pwm_prescale_p1_RNI1QRQ_0_LC_2_14_4.C_ON=1'b0;
    defparam pwm_prescale_p1_RNI1QRQ_0_LC_2_14_4.SEQ_MODE=4'b0000;
    defparam pwm_prescale_p1_RNI1QRQ_0_LC_2_14_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 pwm_prescale_p1_RNI1QRQ_0_LC_2_14_4 (
            .in0(N__4648),
            .in1(N__4596),
            .in2(_gnd_net_),
            .in3(N__4434),
            .lcout(N_38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNO_LC_2_15_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNO_LC_2_15_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNO_LC_2_15_6.LUT_INIT=16'b1000010000100001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_33_c_RNO_LC_2_15_6 (
            .in0(N__3022),
            .in1(N__3001),
            .in2(N__3127),
            .in3(N__3106),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_lout_p1_11_LC_2_16_1.C_ON=1'b0;
    defparam pwm_lout_p1_11_LC_2_16_1.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_11_LC_2_16_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_11_LC_2_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3145),
            .lcout(pwm_lout_p1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4405),
            .ce(),
            .sr(N__4323));
    defparam pwm_lout_p1_10_LC_2_16_6.C_ON=1'b0;
    defparam pwm_lout_p1_10_LC_2_16_6.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_10_LC_2_16_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_10_LC_2_16_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3118),
            .lcout(pwm_lout_p1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4405),
            .ce(),
            .sr(N__4323));
    defparam pwm_lout_p1_1_LC_3_8_2.C_ON=1'b0;
    defparam pwm_lout_p1_1_LC_3_8_2.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_1_LC_3_8_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_1_LC_3_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3100),
            .lcout(pwm_lout_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4397),
            .ce(),
            .sr(N__4319));
    defparam pwm_ctrl_p1_1_LC_3_8_6.C_ON=1'b0;
    defparam pwm_ctrl_p1_1_LC_3_8_6.SEQ_MODE=4'b1010;
    defparam pwm_ctrl_p1_1_LC_3_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_ctrl_p1_1_LC_3_8_6 (
            .in0(N__3085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_ctrl_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4397),
            .ce(),
            .sr(N__4319));
    defparam prescale_cnt_p1_11_LC_3_9_0.C_ON=1'b0;
    defparam prescale_cnt_p1_11_LC_3_9_0.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_11_LC_3_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_11_LC_3_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3772),
            .lcout(prescale_cnt_p1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam pwm_lout_p1_0_LC_3_9_1.C_ON=1'b0;
    defparam pwm_lout_p1_0_LC_3_9_1.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_0_LC_3_9_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_lout_p1_0_LC_3_9_1 (
            .in0(N__3070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_lout_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_cnt_p1_10_LC_3_9_2.C_ON=1'b0;
    defparam prescale_cnt_p1_10_LC_3_9_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_10_LC_3_9_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 prescale_cnt_p1_10_LC_3_9_2 (
            .in0(N__3790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(prescale_cnt_p1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_stop_p1_6_LC_3_9_3.C_ON=1'b0;
    defparam prescale_stop_p1_6_LC_3_9_3.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_6_LC_3_9_3.LUT_INIT=16'b0000010110100000;
    LogicCell40 prescale_stop_p1_6_LC_3_9_3 (
            .in0(N__4491),
            .in1(_gnd_net_),
            .in2(N__4603),
            .in3(N__4667),
            .lcout(prescale_stop_p1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_cnt_p1_7_LC_3_9_4.C_ON=1'b0;
    defparam prescale_cnt_p1_7_LC_3_9_4.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_7_LC_3_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_7_LC_3_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3613),
            .lcout(prescale_cnt_p1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_cnt_p1_6_LC_3_9_5.C_ON=1'b0;
    defparam prescale_cnt_p1_6_LC_3_9_5.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_6_LC_3_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_6_LC_3_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3631),
            .lcout(prescale_cnt_p1Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_stop_p1_10_LC_3_9_6.C_ON=1'b0;
    defparam prescale_stop_p1_10_LC_3_9_6.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_10_LC_3_9_6.LUT_INIT=16'b0010001010001000;
    LogicCell40 prescale_stop_p1_10_LC_3_9_6 (
            .in0(N__4666),
            .in1(N__4599),
            .in2(_gnd_net_),
            .in3(N__4490),
            .lcout(prescale_stop_p1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam prescale_stop_p1_7_LC_3_9_7.C_ON=1'b0;
    defparam prescale_stop_p1_7_LC_3_9_7.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_7_LC_3_9_7.LUT_INIT=16'b0101010100000000;
    LogicCell40 prescale_stop_p1_7_LC_3_9_7 (
            .in0(N__4492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4665),
            .lcout(prescale_stop_p1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4390),
            .ce(),
            .sr(N__4314));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_RNO_LC_3_10_2.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_RNO_LC_3_10_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_RNO_LC_3_10_2.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_39_c_RNO_LC_3_10_2 (
            .in0(N__3301),
            .in1(N__3295),
            .in2(N__3289),
            .in3(N__3280),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_RNO_LC_3_10_3.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_RNO_LC_3_10_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_RNO_LC_3_10_3.LUT_INIT=16'b0010001000010001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_27_c_RNO_LC_3_10_3 (
            .in0(N__3274),
            .in1(N__3268),
            .in2(_gnd_net_),
            .in3(N__3262),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_RNO_LC_3_10_5.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_RNO_LC_3_10_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_1_c_RNO_LC_3_10_5.LUT_INIT=16'b1001000000001001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_1_c_RNO_LC_3_10_5 (
            .in0(N__3255),
            .in1(N__3238),
            .in2(N__3229),
            .in3(N__3208),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctrl_p1_RNI1IE6_0_LC_3_10_6.C_ON=1'b0;
    defparam pwm_ctrl_p1_RNI1IE6_0_LC_3_10_6.SEQ_MODE=4'b0000;
    defparam pwm_ctrl_p1_RNI1IE6_0_LC_3_10_6.LUT_INIT=16'b0000000001010101;
    LogicCell40 pwm_ctrl_p1_RNI1IE6_0_LC_3_10_6 (
            .in0(N__3577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3592),
            .lcout(N_86),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_RNO_LC_3_10_7.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_RNO_LC_3_10_7.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_15_c_RNO_LC_3_10_7.LUT_INIT=16'b1000010000100001;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_15_c_RNO_LC_3_10_7 (
            .in0(N__4003),
            .in1(N__3880),
            .in2(N__3193),
            .in3(N__3170),
            .lcout(proc_pwm_fsm_pwm_loc20_0_N_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_ctrl_p1_RNICQ6G_0_LC_3_11_0.C_ON=1'b0;
    defparam pwm_ctrl_p1_RNICQ6G_0_LC_3_11_0.SEQ_MODE=4'b0000;
    defparam pwm_ctrl_p1_RNICQ6G_0_LC_3_11_0.LUT_INIT=16'b1000100000000000;
    LogicCell40 pwm_ctrl_p1_RNICQ6G_0_LC_3_11_0 (
            .in0(N__3591),
            .in1(N__3576),
            .in2(_gnd_net_),
            .in3(N__3467),
            .lcout(pwm_loc_1_sqmuxa),
            .ltout(pwm_loc_1_sqmuxa_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIMT131_LC_3_11_1.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIMT131_LC_3_11_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIMT131_LC_3_11_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIMT131_LC_3_11_1 (
            .in0(N__3441),
            .in1(_gnd_net_),
            .in2(N__3559),
            .in3(N__3395),
            .lcout(un1_pwm_loc8_1_0),
            .ltout(un1_pwm_loc8_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_tick_RNI46OT1_LC_3_11_2.C_ON=1'b0;
    defparam prescale_tick_RNI46OT1_LC_3_11_2.SEQ_MODE=4'b0000;
    defparam prescale_tick_RNI46OT1_LC_3_11_2.LUT_INIT=16'b1110101011101110;
    LogicCell40 prescale_tick_RNI46OT1_LC_3_11_2 (
            .in0(N__3416),
            .in1(N__3530),
            .in2(N__3556),
            .in3(N__3454),
            .lcout(pwm_cnte_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_togl_LC_3_11_3.C_ON=1'b0;
    defparam pwm_togl_LC_3_11_3.SEQ_MODE=4'b1010;
    defparam pwm_togl_LC_3_11_3.LUT_INIT=16'b0001001000100010;
    LogicCell40 pwm_togl_LC_3_11_3 (
            .in0(N__3443),
            .in1(N__3418),
            .in2(N__3535),
            .in3(N__3541),
            .lcout(pwm_toglZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4391),
            .ce(),
            .sr(N__4305));
    defparam pwm_loc_RNO_1_LC_3_11_4.C_ON=1'b0;
    defparam pwm_loc_RNO_1_LC_3_11_4.SEQ_MODE=4'b0000;
    defparam pwm_loc_RNO_1_LC_3_11_4.LUT_INIT=16'b1100010000000100;
    LogicCell40 pwm_loc_RNO_1_LC_3_11_4 (
            .in0(N__3397),
            .in1(N__3529),
            .in2(N__3448),
            .in3(N__3505),
            .lcout(),
            .ltout(pwm_loc_1_sqmuxa_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwm_loc_LC_3_11_5.C_ON=1'b0;
    defparam pwm_loc_LC_3_11_5.SEQ_MODE=4'b1010;
    defparam pwm_loc_LC_3_11_5.LUT_INIT=16'b1100110001010100;
    LogicCell40 pwm_loc_LC_3_11_5 (
            .in0(N__3499),
            .in1(N__3480),
            .in2(N__3493),
            .in3(N__3417),
            .lcout(pwm_locZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4391),
            .ce(),
            .sr(N__4305));
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNIKR9E_LC_3_11_6.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNIKR9E_LC_3_11_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc20_0_I_33_c_RNIKR9E_LC_3_11_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 proc_pwm_fsm_pwm_loc20_0_I_33_c_RNIKR9E_LC_3_11_6 (
            .in0(_gnd_net_),
            .in1(N__3440),
            .in2(_gnd_net_),
            .in3(N__3468),
            .lcout(N_87),
            .ltout(N_87_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIVGJ71_LC_3_11_7.C_ON=1'b0;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIVGJ71_LC_3_11_7.SEQ_MODE=4'b0000;
    defparam proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIVGJ71_LC_3_11_7.LUT_INIT=16'b1111110111111100;
    LogicCell40 proc_pwm_fsm_pwm_loc8_0_I_33_c_RNIVGJ71_LC_3_11_7 (
            .in0(N__3442),
            .in1(N__3415),
            .in2(N__3400),
            .in3(N__3396),
            .lcout(N_78_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_RNO_0_0_LC_3_12_0.C_ON=1'b1;
    defparam prescale_cnt_RNO_0_0_LC_3_12_0.SEQ_MODE=4'b0000;
    defparam prescale_cnt_RNO_0_0_LC_3_12_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 prescale_cnt_RNO_0_0_LC_3_12_0 (
            .in0(_gnd_net_),
            .in1(N__3321),
            .in2(_gnd_net_),
            .in3(N__3304),
            .lcout(prescale_cnt_s_0),
            .ltout(),
            .carryin(bfn_3_12_0_),
            .carryout(prescale_cnt_cry_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_1_LC_3_12_1.C_ON=1'b1;
    defparam prescale_cnt_1_LC_3_12_1.SEQ_MODE=4'b1010;
    defparam prescale_cnt_1_LC_3_12_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_1_LC_3_12_1 (
            .in0(N__3738),
            .in1(N__3657),
            .in2(_gnd_net_),
            .in3(N__3646),
            .lcout(prescale_cntZ0Z_1),
            .ltout(),
            .carryin(prescale_cnt_cry_0),
            .carryout(prescale_cnt_cry_1),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_2_LC_3_12_2.C_ON=1'b1;
    defparam prescale_cnt_2_LC_3_12_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_2_LC_3_12_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_2_LC_3_12_2 (
            .in0(N__3731),
            .in1(N__4125),
            .in2(_gnd_net_),
            .in3(N__3643),
            .lcout(prescale_cntZ0Z_2),
            .ltout(),
            .carryin(prescale_cnt_cry_1),
            .carryout(prescale_cnt_cry_2),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_3_LC_3_12_3.C_ON=1'b1;
    defparam prescale_cnt_3_LC_3_12_3.SEQ_MODE=4'b1010;
    defparam prescale_cnt_3_LC_3_12_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_3_LC_3_12_3 (
            .in0(N__3739),
            .in1(N__4149),
            .in2(_gnd_net_),
            .in3(N__3640),
            .lcout(prescale_cntZ0Z_3),
            .ltout(),
            .carryin(prescale_cnt_cry_2),
            .carryout(prescale_cnt_cry_3),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_4_LC_3_12_4.C_ON=1'b1;
    defparam prescale_cnt_4_LC_3_12_4.SEQ_MODE=4'b1010;
    defparam prescale_cnt_4_LC_3_12_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_4_LC_3_12_4 (
            .in0(N__3732),
            .in1(N__4716),
            .in2(_gnd_net_),
            .in3(N__3637),
            .lcout(prescale_cntZ0Z_4),
            .ltout(),
            .carryin(prescale_cnt_cry_3),
            .carryout(prescale_cnt_cry_4),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_5_LC_3_12_5.C_ON=1'b1;
    defparam prescale_cnt_5_LC_3_12_5.SEQ_MODE=4'b1010;
    defparam prescale_cnt_5_LC_3_12_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_5_LC_3_12_5 (
            .in0(N__3740),
            .in1(N__3864),
            .in2(_gnd_net_),
            .in3(N__3634),
            .lcout(prescale_cntZ0Z_5),
            .ltout(),
            .carryin(prescale_cnt_cry_4),
            .carryout(prescale_cnt_cry_5),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_6_LC_3_12_6.C_ON=1'b1;
    defparam prescale_cnt_6_LC_3_12_6.SEQ_MODE=4'b1010;
    defparam prescale_cnt_6_LC_3_12_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_6_LC_3_12_6 (
            .in0(N__3733),
            .in1(N__3627),
            .in2(_gnd_net_),
            .in3(N__3616),
            .lcout(prescale_cntZ0Z_6),
            .ltout(),
            .carryin(prescale_cnt_cry_5),
            .carryout(prescale_cnt_cry_6),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_7_LC_3_12_7.C_ON=1'b1;
    defparam prescale_cnt_7_LC_3_12_7.SEQ_MODE=4'b1010;
    defparam prescale_cnt_7_LC_3_12_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_7_LC_3_12_7 (
            .in0(N__3741),
            .in1(N__3609),
            .in2(_gnd_net_),
            .in3(N__3598),
            .lcout(prescale_cntZ0Z_7),
            .ltout(),
            .carryin(prescale_cnt_cry_6),
            .carryout(prescale_cnt_cry_7),
            .clk(N__4398),
            .ce(),
            .sr(N__4311));
    defparam prescale_cnt_8_LC_3_13_0.C_ON=1'b1;
    defparam prescale_cnt_8_LC_3_13_0.SEQ_MODE=4'b1010;
    defparam prescale_cnt_8_LC_3_13_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_8_LC_3_13_0 (
            .in0(N__3730),
            .in1(N__3978),
            .in2(_gnd_net_),
            .in3(N__3595),
            .lcout(prescale_cntZ0Z_8),
            .ltout(),
            .carryin(bfn_3_13_0_),
            .carryout(prescale_cnt_cry_8),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_9_LC_3_13_1.C_ON=1'b1;
    defparam prescale_cnt_9_LC_3_13_1.SEQ_MODE=4'b1010;
    defparam prescale_cnt_9_LC_3_13_1.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_9_LC_3_13_1 (
            .in0(N__3737),
            .in1(N__3954),
            .in2(_gnd_net_),
            .in3(N__3793),
            .lcout(prescale_cntZ0Z_9),
            .ltout(),
            .carryin(prescale_cnt_cry_8),
            .carryout(prescale_cnt_cry_9),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_10_LC_3_13_2.C_ON=1'b1;
    defparam prescale_cnt_10_LC_3_13_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_10_LC_3_13_2.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_10_LC_3_13_2 (
            .in0(N__3727),
            .in1(N__3786),
            .in2(_gnd_net_),
            .in3(N__3775),
            .lcout(prescale_cntZ0Z_10),
            .ltout(),
            .carryin(prescale_cnt_cry_9),
            .carryout(prescale_cnt_cry_10),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_11_LC_3_13_3.C_ON=1'b1;
    defparam prescale_cnt_11_LC_3_13_3.SEQ_MODE=4'b1010;
    defparam prescale_cnt_11_LC_3_13_3.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_11_LC_3_13_3 (
            .in0(N__3734),
            .in1(N__3768),
            .in2(_gnd_net_),
            .in3(N__3757),
            .lcout(prescale_cntZ0Z_11),
            .ltout(),
            .carryin(prescale_cnt_cry_10),
            .carryout(prescale_cnt_cry_11),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_12_LC_3_13_4.C_ON=1'b1;
    defparam prescale_cnt_12_LC_3_13_4.SEQ_MODE=4'b1010;
    defparam prescale_cnt_12_LC_3_13_4.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_12_LC_3_13_4 (
            .in0(N__3728),
            .in1(N__4203),
            .in2(_gnd_net_),
            .in3(N__3754),
            .lcout(prescale_cntZ0Z_12),
            .ltout(),
            .carryin(prescale_cnt_cry_11),
            .carryout(prescale_cnt_cry_12),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_13_LC_3_13_5.C_ON=1'b1;
    defparam prescale_cnt_13_LC_3_13_5.SEQ_MODE=4'b1010;
    defparam prescale_cnt_13_LC_3_13_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_13_LC_3_13_5 (
            .in0(N__3735),
            .in1(N__4101),
            .in2(_gnd_net_),
            .in3(N__3751),
            .lcout(prescale_cntZ0Z_13),
            .ltout(),
            .carryin(prescale_cnt_cry_12),
            .carryout(prescale_cnt_cry_13),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_14_LC_3_13_6.C_ON=1'b1;
    defparam prescale_cnt_14_LC_3_13_6.SEQ_MODE=4'b1010;
    defparam prescale_cnt_14_LC_3_13_6.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_14_LC_3_13_6 (
            .in0(N__3729),
            .in1(N__3837),
            .in2(_gnd_net_),
            .in3(N__3748),
            .lcout(prescale_cntZ0Z_14),
            .ltout(),
            .carryin(prescale_cnt_cry_13),
            .carryout(prescale_cnt_cry_14),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_15_LC_3_13_7.C_ON=1'b1;
    defparam prescale_cnt_15_LC_3_13_7.SEQ_MODE=4'b1010;
    defparam prescale_cnt_15_LC_3_13_7.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_15_LC_3_13_7 (
            .in0(N__3736),
            .in1(N__3810),
            .in2(_gnd_net_),
            .in3(N__3745),
            .lcout(prescale_cntZ0Z_15),
            .ltout(),
            .carryin(prescale_cnt_cry_14),
            .carryout(prescale_cnt_cry_15),
            .clk(N__4399),
            .ce(),
            .sr(N__4315));
    defparam prescale_cnt_16_LC_3_14_0.C_ON=1'b0;
    defparam prescale_cnt_16_LC_3_14_0.SEQ_MODE=4'b1010;
    defparam prescale_cnt_16_LC_3_14_0.LUT_INIT=16'b0001000101000100;
    LogicCell40 prescale_cnt_16_LC_3_14_0 (
            .in0(N__3742),
            .in1(N__4188),
            .in2(_gnd_net_),
            .in3(N__3679),
            .lcout(prescale_cntZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4403),
            .ce(),
            .sr(N__4320));
    defparam prescale_stop_p1_0_LC_3_14_6.C_ON=1'b0;
    defparam prescale_stop_p1_0_LC_3_14_6.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_0_LC_3_14_6.LUT_INIT=16'b1111111111101110;
    LogicCell40 prescale_stop_p1_0_LC_3_14_6 (
            .in0(N__4678),
            .in1(N__4597),
            .in2(_gnd_net_),
            .in3(N__4461),
            .lcout(prescale_stop_p1Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4403),
            .ce(),
            .sr(N__4320));
    defparam prescale_stop_p1_1_LC_3_14_7.C_ON=1'b0;
    defparam prescale_stop_p1_1_LC_3_14_7.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_1_LC_3_14_7.LUT_INIT=16'b1111111110001000;
    LogicCell40 prescale_stop_p1_1_LC_3_14_7 (
            .in0(N__4462),
            .in1(N__4598),
            .in2(_gnd_net_),
            .in3(N__4679),
            .lcout(prescale_stop_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4403),
            .ce(),
            .sr(N__4320));
    defparam pwm_lout_p1_4_LC_3_18_3.C_ON=1'b0;
    defparam pwm_lout_p1_4_LC_3_18_3.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_4_LC_3_18_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_4_LC_3_18_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3898),
            .lcout(pwm_lout_p1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4408),
            .ce(),
            .sr(N__4327));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_RNO_LC_5_8_0.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_RNO_LC_5_8_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_RNO_LC_5_8_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_15_c_RNO_LC_5_8_0 (
            .in0(N__4227),
            .in1(N__3799),
            .in2(N__3853),
            .in3(N__3826),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_p1_5_LC_5_9_0.C_ON=1'b0;
    defparam prescale_cnt_p1_5_LC_5_9_0.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_5_LC_5_9_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_5_LC_5_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3871),
            .lcout(prescale_cnt_p1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4400),
            .ce(),
            .sr(N__4324));
    defparam prescale_stop_p1_14_LC_5_9_1.C_ON=1'b0;
    defparam prescale_stop_p1_14_LC_5_9_1.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_14_LC_5_9_1.LUT_INIT=16'b1000100000000000;
    LogicCell40 prescale_stop_p1_14_LC_5_9_1 (
            .in0(N__4687),
            .in1(N__4573),
            .in2(_gnd_net_),
            .in3(N__4489),
            .lcout(prescale_stop_p1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4400),
            .ce(),
            .sr(N__4324));
    defparam prescale_stop_p1_15_LC_5_9_4.C_ON=1'b0;
    defparam prescale_stop_p1_15_LC_5_9_4.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_15_LC_5_9_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 prescale_stop_p1_15_LC_5_9_4 (
            .in0(N__4574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4162),
            .lcout(prescale_stop_p1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4400),
            .ce(),
            .sr(N__4324));
    defparam prescale_cnt_p1_14_LC_5_9_6.C_ON=1'b0;
    defparam prescale_cnt_p1_14_LC_5_9_6.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_14_LC_5_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_14_LC_5_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3844),
            .lcout(prescale_cnt_p1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4400),
            .ce(),
            .sr(N__4324));
    defparam prescale_cnt_p1_15_LC_5_9_7.C_ON=1'b0;
    defparam prescale_cnt_p1_15_LC_5_9_7.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_15_LC_5_9_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_15_LC_5_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3820),
            .lcout(prescale_cnt_p1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4400),
            .ce(),
            .sr(N__4324));
    defparam prescale_stop_p1_8_LC_5_10_1.C_ON=1'b0;
    defparam prescale_stop_p1_8_LC_5_10_1.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_8_LC_5_10_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 prescale_stop_p1_8_LC_5_10_1 (
            .in0(_gnd_net_),
            .in1(N__4688),
            .in2(_gnd_net_),
            .in3(N__4572),
            .lcout(prescale_stop_p1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4392),
            .ce(),
            .sr(N__4321));
    defparam prescale_stop_p1_2_LC_5_10_3.C_ON=1'b0;
    defparam prescale_stop_p1_2_LC_5_10_3.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_2_LC_5_10_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_stop_p1_2_LC_5_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4689),
            .lcout(prescale_stop_p1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4392),
            .ce(),
            .sr(N__4321));
    defparam pwm_prescale_p1_1_LC_5_10_4.C_ON=1'b0;
    defparam pwm_prescale_p1_1_LC_5_10_4.SEQ_MODE=4'b1010;
    defparam pwm_prescale_p1_1_LC_5_10_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 pwm_prescale_p1_1_LC_5_10_4 (
            .in0(N__4030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pwm_prescale_p1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4392),
            .ce(),
            .sr(N__4321));
    defparam pwm_lout_p1_5_LC_5_10_7.C_ON=1'b0;
    defparam pwm_lout_p1_5_LC_5_10_7.SEQ_MODE=4'b1010;
    defparam pwm_lout_p1_5_LC_5_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 pwm_lout_p1_5_LC_5_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4021),
            .lcout(pwm_lout_p1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4392),
            .ce(),
            .sr(N__4321));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_RNO_LC_5_11_0.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_RNO_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_RNO_LC_5_11_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_33_c_RNO_LC_5_11_0 (
            .in0(N__3943),
            .in1(N__3967),
            .in2(N__3994),
            .in3(N__3937),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_p1_8_LC_5_11_1.C_ON=1'b0;
    defparam prescale_cnt_p1_8_LC_5_11_1.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_8_LC_5_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_8_LC_5_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3985),
            .lcout(prescale_cnt_p1Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4401),
            .ce(),
            .sr(N__4312));
    defparam prescale_cnt_p1_9_LC_5_11_2.C_ON=1'b0;
    defparam prescale_cnt_p1_9_LC_5_11_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_9_LC_5_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_9_LC_5_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3961),
            .lcout(prescale_cnt_p1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4401),
            .ce(),
            .sr(N__4312));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_RNO_LC_5_11_5.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_RNO_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_RNO_LC_5_11_5.LUT_INIT=16'b1000001001000001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_51_c_RNO_LC_5_11_5 (
            .in0(N__3936),
            .in1(N__4138),
            .in2(N__3928),
            .in3(N__4114),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_stop_p1_3_LC_5_11_7.C_ON=1'b0;
    defparam prescale_stop_p1_3_LC_5_11_7.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_3_LC_5_11_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 prescale_stop_p1_3_LC_5_11_7 (
            .in0(N__4698),
            .in1(N__4575),
            .in2(_gnd_net_),
            .in3(N__4478),
            .lcout(prescale_stop_p1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4401),
            .ce(),
            .sr(N__4312));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_LC_5_12_0.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_LC_5_12_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_1_c_LC_5_12_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_1_c_LC_5_12_0 (
            .in0(_gnd_net_),
            .in1(N__3919),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_12_0_),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_0),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_LC_5_12_1.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_51_c_LC_5_12_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_51_c_LC_5_12_1 (
            .in0(_gnd_net_),
            .in1(N__4090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_0),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_LC_5_12_2.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_LC_5_12_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_45_c_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__4237),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_1),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_LC_5_12_3.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_LC_5_12_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_39_c_LC_5_12_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_39_c_LC_5_12_3 (
            .in0(_gnd_net_),
            .in1(N__4084),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_2),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_LC_5_12_4.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_LC_5_12_4.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_33_c_LC_5_12_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_33_c_LC_5_12_4 (
            .in0(_gnd_net_),
            .in1(N__4072),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_3),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_LC_5_12_5.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_LC_5_12_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_27_c_LC_5_12_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_27_c_LC_5_12_5 (
            .in0(_gnd_net_),
            .in1(N__4066),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_4),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_LC_5_12_6.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_LC_5_12_6.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_LC_5_12_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_21_c_LC_5_12_6 (
            .in0(_gnd_net_),
            .in1(N__4504),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_5),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_LC_5_12_7.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_LC_5_12_7.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_15_c_LC_5_12_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_15_c_LC_5_12_7 (
            .in0(_gnd_net_),
            .in1(N__4054),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(proc_pwm_cnt_prescale_cnt10_0_data_tmp_6),
            .carryout(proc_pwm_cnt_prescale_cnt10_0_data_tmp_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_LC_5_13_0.C_ON=1'b1;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_LC_5_13_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_9_c_LC_5_13_0 (
            .in0(_gnd_net_),
            .in1(N__4216),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(proc_pwm_cnt_prescale_cnt10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_THRU_LUT4_0_LC_5_13_1.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_THRU_LUT4_0_LC_5_13_1.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_THRU_LUT4_0_LC_5_13_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_THRU_LUT4_0_LC_5_13_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4045),
            .lcout(proc_pwm_cnt_prescale_cnt10_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_RNO_LC_5_13_2.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_RNO_LC_5_13_2.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_45_c_RNO_LC_5_13_2.LUT_INIT=16'b1001000000001001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_45_c_RNO_LC_5_13_2 (
            .in0(N__4728),
            .in1(N__4705),
            .in2(N__4171),
            .in3(N__4246),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNO_LC_5_13_3.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNO_LC_5_13_3.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNO_LC_5_13_3.LUT_INIT=16'b0000000010011001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_9_c_RNO_LC_5_13_3 (
            .in0(N__4177),
            .in1(N__4729),
            .in2(_gnd_net_),
            .in3(N__4231),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_36),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_p1_12_LC_5_14_0.C_ON=1'b0;
    defparam prescale_cnt_p1_12_LC_5_14_0.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_12_LC_5_14_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_12_LC_5_14_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4210),
            .lcout(prescale_cnt_p1Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4406),
            .ce(),
            .sr(N__4325));
    defparam prescale_cnt_p1_16_LC_5_14_2.C_ON=1'b0;
    defparam prescale_cnt_p1_16_LC_5_14_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_16_LC_5_14_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 prescale_cnt_p1_16_LC_5_14_2 (
            .in0(N__4192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(prescale_cnt_p1Z0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4406),
            .ce(),
            .sr(N__4325));
    defparam prescale_stop_p1_5_LC_5_14_4.C_ON=1'b0;
    defparam prescale_stop_p1_5_LC_5_14_4.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_5_LC_5_14_4.LUT_INIT=16'b1100110000100010;
    LogicCell40 prescale_stop_p1_5_LC_5_14_4 (
            .in0(N__4699),
            .in1(N__4595),
            .in2(_gnd_net_),
            .in3(N__4479),
            .lcout(prescale_stop_p1Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4406),
            .ce(),
            .sr(N__4325));
    defparam prescale_stop_1_8_3__m8_0_a3_LC_6_9_4.C_ON=1'b0;
    defparam prescale_stop_1_8_3__m8_0_a3_LC_6_9_4.SEQ_MODE=4'b0000;
    defparam prescale_stop_1_8_3__m8_0_a3_LC_6_9_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 prescale_stop_1_8_3__m8_0_a3_LC_6_9_4 (
            .in0(_gnd_net_),
            .in1(N__4680),
            .in2(_gnd_net_),
            .in3(N__4488),
            .lcout(prescale_stop_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_cnt_p1_3_LC_6_11_2.C_ON=1'b0;
    defparam prescale_cnt_p1_3_LC_6_11_2.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_3_LC_6_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_3_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4156),
            .lcout(prescale_cnt_p1Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4402),
            .ce(),
            .sr(N__4316));
    defparam prescale_cnt_p1_2_LC_6_11_6.C_ON=1'b0;
    defparam prescale_cnt_p1_2_LC_6_11_6.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_2_LC_6_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_2_LC_6_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4132),
            .lcout(prescale_cnt_p1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4402),
            .ce(),
            .sr(N__4316));
    defparam prescale_cnt_p1_13_LC_6_11_7.C_ON=1'b0;
    defparam prescale_cnt_p1_13_LC_6_11_7.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_13_LC_6_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_13_LC_6_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4108),
            .lcout(prescale_cnt_p1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4402),
            .ce(),
            .sr(N__4316));
    defparam prescale_stop_p1_4_LC_6_12_0.C_ON=1'b0;
    defparam prescale_stop_p1_4_LC_6_12_0.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_4_LC_6_12_0.LUT_INIT=16'b1100110000000000;
    LogicCell40 prescale_stop_p1_4_LC_6_12_0 (
            .in0(_gnd_net_),
            .in1(N__4594),
            .in2(_gnd_net_),
            .in3(N__4697),
            .lcout(prescale_stop_p1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4404),
            .ce(),
            .sr(N__4322));
    defparam prescale_cnt_p1_4_LC_6_12_1.C_ON=1'b0;
    defparam prescale_cnt_p1_4_LC_6_12_1.SEQ_MODE=4'b1010;
    defparam prescale_cnt_p1_4_LC_6_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 prescale_cnt_p1_4_LC_6_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4720),
            .lcout(prescale_cnt_p1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4404),
            .ce(),
            .sr(N__4322));
    defparam prescale_stop_1_8_3__m4_0_a3_LC_6_13_2.C_ON=1'b0;
    defparam prescale_stop_1_8_3__m4_0_a3_LC_6_13_2.SEQ_MODE=4'b0000;
    defparam prescale_stop_1_8_3__m4_0_a3_LC_6_13_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 prescale_stop_1_8_3__m4_0_a3_LC_6_13_2 (
            .in0(_gnd_net_),
            .in1(N__4696),
            .in2(_gnd_net_),
            .in3(N__4593),
            .lcout(prescale_stop_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_RNO_LC_6_13_5.C_ON=1'b0;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_RNO_LC_6_13_5.SEQ_MODE=4'b0000;
    defparam proc_pwm_cnt_prescale_cnt10_0_I_21_c_RNO_LC_6_13_5.LUT_INIT=16'b0000000010011001;
    LogicCell40 proc_pwm_cnt_prescale_cnt10_0_I_21_c_RNO_LC_6_13_5 (
            .in0(N__4414),
            .in1(N__4519),
            .in2(_gnd_net_),
            .in3(N__4510),
            .lcout(proc_pwm_cnt_prescale_cnt10_0_N_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam prescale_stop_p1_13_LC_6_14_2.C_ON=1'b0;
    defparam prescale_stop_p1_13_LC_6_14_2.SEQ_MODE=4'b1010;
    defparam prescale_stop_p1_13_LC_6_14_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 prescale_stop_p1_13_LC_6_14_2 (
            .in0(_gnd_net_),
            .in1(N__4498),
            .in2(_gnd_net_),
            .in3(N__4480),
            .lcout(prescale_stop_p1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4407),
            .ce(),
            .sr(N__4326));
endmodule // gpio_pwm
